// SPDX-License-Identifier: GPL-3.0-only
/*
 * GW2AR-LV18QN88C8/I7 SDRAM controller
 *
 * Copyright (C) 2023 Luís Mendes <luis.p.mendes@gmail.com>
 */
/* PageWords= 256, Address width: 8 *)
/* Number of Read/Write suspend cycles/wait states    : 0 *)
/* Row cycle time (same bank)                   - RC  : 7 */
/* RAS to CAS delay (same bank)                 - RCD : 6 */
/* PreCharge to Refresh/Row activate (same bank)- RP  : 2 */
/* Row activate to row activate (diff. banks)   - RRD : 2 */
/* Row activate to pre-charge cycles (same bank)- RAS : 5 */
/* Write recovery time                          - WR  : 2 */
/* Mode register set cycle cycles               - MRD : 4 */
/* Average refresh interval cycles              - REFI: 936 */
/* Mask bit offset                                    : 0 */
/* Column address width                               : 8 */
/* Bank address width                                 : 2 */
/* Row address width                                  : 11 */
/* Generated by Yosys 0.17+9 (git sha1 98c7804b8, clang 10.0.0-4ubuntu1 -fPIC -Os) */

(* \amaranth.hierarchy  = "top.sdramController.bankController0" *)
(* generator = "Amaranth" *)
module bankController0(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$1  = 0;
  (* src = "sdram_controller.py:1189" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1190" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1212" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1217" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1177" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1175" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1169" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1169" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1174" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1178" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1172" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1172" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1189" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1190" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1189" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1189" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1192" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1198" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$36  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1198" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1201" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1208" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1208" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1208" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1212" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1213" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1217" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1189" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1218" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1190" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1190" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1199" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1202" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* src = "sdram_controller.py:1199" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1210" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1210" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h6;
      /* src = "sdram_controller.py:1212" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1215" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1215" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1217" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController.bankController1" *)
(* generator = "Amaranth" *)
module bankController1(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$2  = 0;
  (* src = "sdram_controller.py:1189" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1190" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1212" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1217" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1177" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1175" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1169" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1169" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1174" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1178" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1172" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1172" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1189" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1190" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1189" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1189" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1192" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1198" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$36  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1198" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1201" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1208" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1208" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1208" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1212" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1213" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1217" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1189" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1218" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1190" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1190" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1199" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1202" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* src = "sdram_controller.py:1199" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1210" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1210" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h6;
      /* src = "sdram_controller.py:1212" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1215" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1215" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1217" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController.bankController2" *)
(* generator = "Amaranth" *)
module bankController2(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$3  = 0;
  (* src = "sdram_controller.py:1189" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1190" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1212" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1217" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1177" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1175" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1169" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1169" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1174" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1178" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1172" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1172" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1189" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1190" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1189" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1189" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1192" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1198" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$36  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1198" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1201" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1208" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1208" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1208" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1212" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1213" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1217" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1189" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1218" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1190" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1190" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1199" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1202" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* src = "sdram_controller.py:1199" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1210" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1210" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h6;
      /* src = "sdram_controller.py:1212" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1215" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1215" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1217" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController.bankController3" *)
(* generator = "Amaranth" *)
module bankController3(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$4  = 0;
  (* src = "sdram_controller.py:1189" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1190" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1191" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1198" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1199" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1201" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1208" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1212" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1213" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1217" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1218" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1189" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1177" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1171" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1175" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1170" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1169" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1169" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1174" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1288" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1178" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1172" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1172" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1189" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1190" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1189" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1189" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1189" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1192" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1198" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$36  = bankState == (* src = "sdram_controller.py:1198" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1198" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1189" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1198" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1199" *) 3'h4;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1201" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1208" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1208" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1208" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1212" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1213" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1217" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1189" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1218" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1189" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1190" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1190" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1189" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1189" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1194" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1199" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1202" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1198" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1198" */
      1'h1:
          (* src = "sdram_controller.py:1199" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1199" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1204" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1210" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1210" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h6;
      /* src = "sdram_controller.py:1212" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1215" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1215" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1217" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController" *)
(* generator = "Amaranth" *)
module sdramController(sdramClkEn, sdramCSn, sdramRASn, sdramCASn, sdramWEn, sdramAddress, sdramBank, ctrlReady, ctrlRd, ctrlWr, ctrlRdAddress, ctrlWrAddress, sdramDataMasks, ctrlRdIncAddress, ctrlRdDataOut, sdramDqOut, ctrlWrIncAddress, sdramDqWRn, sdramDqIn, ctrlWrDataIn, sdramClk
);
  reg \$auto$verilog_backend.cc:2083:dump_module$5  = 0;
  (* src = "sdram_controller.py:655" *)
  wire \$1 ;
  (* src = "sdram_controller.py:712" *)
  wire \$1000 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1002 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1004 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1006 ;
  (* src = "sdram_controller.py:483" *)
  wire \$1008 ;
  (* src = "sdram_controller.py:970" *)
  wire \$101 ;
  (* src = "sdram_controller.py:489" *)
  wire \$1010 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1012 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1014 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1016 ;
  (* src = "sdram_controller.py:508" *)
  wire \$1018 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1020 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1022 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1024 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1026 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1028 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$103 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1030 ;
  (* src = "sdram_controller.py:837" *)
  wire \$1032 ;
  (* src = "sdram_controller.py:838" *)
  wire \$1034 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1036 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1038 ;
  (* src = "sdram_controller.py:440" *)
  wire \$1040 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1042 ;
  (* src = "sdram_controller.py:446" *)
  wire \$1044 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1046 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1048 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$105 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1050 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1052 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1054 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1056 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1058 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1060 ;
  (* src = "sdram_controller.py:965" *)
  wire \$1062 ;
  (* src = "sdram_controller.py:508" *)
  wire \$1064 ;
  (* src = "sdram_controller.py:970" *)
  wire \$1066 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$1068 ;
  (* src = "sdram_controller.py:1020" *)
  wire \$107 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1070 ;
  (* src = "sdram_controller.py:396" *)
  wire \$1072 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1074 ;
  (* src = "sdram_controller.py:402" *)
  wire \$1076 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1078 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1080 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1082 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1084 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1086 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1088 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$109 ;
  (* src = "sdram_controller.py:712" *)
  wire \$1090 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1092 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1094 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1096 ;
  (* src = "sdram_controller.py:483" *)
  wire \$1098 ;
  (* src = "sdram_controller.py:723" *)
  wire \$11 ;
  (* src = "sdram_controller.py:489" *)
  wire \$1100 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1102 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1104 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1106 ;
  (* src = "sdram_controller.py:508" *)
  wire \$1108 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$111 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1110 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1112 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1114 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1116 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1118 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1120 ;
  (* src = "sdram_controller.py:837" *)
  wire \$1122 ;
  (* src = "sdram_controller.py:838" *)
  wire \$1124 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1126 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1128 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$113 ;
  (* src = "sdram_controller.py:440" *)
  wire \$1130 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1132 ;
  (* src = "sdram_controller.py:446" *)
  wire \$1134 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1136 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1138 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1140 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1142 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1144 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1146 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1148 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$115 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1150 ;
  (* src = "sdram_controller.py:965" *)
  wire \$1152 ;
  (* src = "sdram_controller.py:508" *)
  wire \$1154 ;
  (* src = "sdram_controller.py:970" *)
  wire \$1156 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$1158 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1160 ;
  (* src = "sdram_controller.py:396" *)
  wire \$1162 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1164 ;
  (* src = "sdram_controller.py:402" *)
  wire \$1166 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1168 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$117 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1170 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1172 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1174 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1176 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1178 ;
  (* src = "sdram_controller.py:722" *)
  wire \$1180 ;
  (* src = "sdram_controller.py:723" *)
  wire \$1182 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1184 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1186 ;
  (* src = "sdram_controller.py:386" *)
  wire \$1188 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$119 ;
  (* src = "sdram_controller.py:388" *)
  wire \$1190 ;
  (* src = "sdram_controller.py:387" *)
  wire [4:0] \$1192 ;
  (* src = "sdram_controller.py:387" *)
  wire [4:0] \$1193 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1195 ;
  (* src = "sdram_controller.py:483" *)
  wire \$1197 ;
  (* src = "sdram_controller.py:489" *)
  wire \$1199 ;
  (* src = "sdram_controller.py:497" *)
  wire \$1201 ;
  (* src = "sdram_controller.py:499" *)
  wire \$1203 ;
  (* src = "sdram_controller.py:498" *)
  wire [4:0] \$1205 ;
  (* src = "sdram_controller.py:498" *)
  wire [4:0] \$1206 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1208 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$121 ;
  (* src = "sdram_controller.py:763" *)
  wire \$1210 ;
  (* src = "sdram_controller.py:764" *)
  wire \$1212 ;
  (* src = "sdram_controller.py:766" *)
  wire \$1214 ;
  (* src = "sdram_controller.py:765" *)
  wire [4:0] \$1216 ;
  (* src = "sdram_controller.py:765" *)
  wire [4:0] \$1217 ;
  (* src = "sdram_controller.py:831" *)
  wire \$1219 ;
  (* src = "sdram_controller.py:837" *)
  wire \$1221 ;
  (* src = "sdram_controller.py:838" *)
  wire \$1223 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1225 ;
  (* src = "sdram_controller.py:839" *)
  wire [4:0] \$1227 ;
  (* src = "sdram_controller.py:839" *)
  wire [4:0] \$1228 ;
  (* src = "sdram_controller.py:712" *)
  wire \$123 ;
  (* src = "sdram_controller.py:926" *)
  wire \$1230 ;
  (* src = "sdram_controller.py:932" *)
  wire \$1232 ;
  (* src = "sdram_controller.py:934" *)
  wire \$1234 ;
  (* src = "sdram_controller.py:935" *)
  wire [4:0] \$1236 ;
  (* src = "sdram_controller.py:935" *)
  wire [4:0] \$1237 ;
  (* src = "sdram_controller.py:936" *)
  wire \$1239 ;
  (* src = "sdram_controller.py:965" *)
  wire \$1241 ;
  (* src = "sdram_controller.py:970" *)
  wire \$1243 ;
  (* src = "sdram_controller.py:997" *)
  wire \$1245 ;
  (* src = "sdram_controller.py:998" *)
  wire [4:0] \$1247 ;
  (* src = "sdram_controller.py:998" *)
  wire [4:0] \$1248 ;
  (* src = "sdram_controller.py:737" *)
  wire \$125 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$1250 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$1252 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$1254 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$1256 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$1258 ;
  (* src = "sdram_controller.py:1066" *)
  wire [4:0] \$1260 ;
  (* src = "sdram_controller.py:1066" *)
  wire [4:0] \$1261 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1263 ;
  (* src = "sdram_controller.py:1070" *)
  wire \$1265 ;
  (* src = "sdram_controller.py:1071" *)
  wire [4:0] \$1267 ;
  (* src = "sdram_controller.py:1071" *)
  wire [4:0] \$1268 ;
  (* src = "sdram_controller.py:742" *)
  wire \$127 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1270 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$1272 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$1274 ;
  (* src = "sdram_controller.py:1081" *)
  wire [4:0] \$1276 ;
  (* src = "sdram_controller.py:1081" *)
  wire [4:0] \$1277 ;
  (* src = "sdram_controller.py:1082" *)
  wire \$1279 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1281 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$1283 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1285 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1287 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1289 ;
  (* src = "sdram_controller.py:746" *)
  wire \$129 ;
  (* src = "sdram_controller.py:1102" *)
  wire [4:0] \$1291 ;
  (* src = "sdram_controller.py:1102" *)
  wire [4:0] \$1292 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1294 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1296 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1298 ;
  (* src = "sdram_controller.py:769" *)
  wire \$13 ;
  (* src = "sdram_controller.py:748" *)
  wire \$1300 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1302 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1304 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1306 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1308 ;
  (* src = "sdram_controller.py:754" *)
  wire \$131 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1310 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1312 ;
  (* src = "sdram_controller.py:837" *)
  wire \$1314 ;
  (* src = "sdram_controller.py:838" *)
  wire \$1316 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1318 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1320 ;
  (* src = "sdram_controller.py:440" *)
  wire \$1322 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1324 ;
  (* src = "sdram_controller.py:446" *)
  wire \$1326 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1328 ;
  (* src = "sdram_controller.py:758" *)
  wire \$133 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1330 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1332 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1334 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1336 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1338 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1340 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1342 ;
  (* src = "sdram_controller.py:970" *)
  wire \$1344 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$1346 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1348 ;
  (* src = "sdram_controller.py:820" *)
  wire \$135 ;
  (* src = "sdram_controller.py:396" *)
  wire \$1350 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1352 ;
  (* src = "sdram_controller.py:402" *)
  wire \$1354 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1356 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1358 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1360 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1362 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1364 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1366 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1368 ;
  (* src = "sdram_controller.py:831" *)
  wire \$137 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1370 ;
  (* src = "sdram_controller.py:769" *)
  wire \$1372 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1374 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1376 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1378 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1380 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1382 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1384 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1386 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1388 ;
  (* src = "sdram_controller.py:837" *)
  wire \$139 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1390 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1392 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1394 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1396 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1398 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1400 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1402 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1404 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1406 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1408 ;
  (* src = "sdram_controller.py:838" *)
  wire \$141 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1410 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1412 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1414 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1416 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1418 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1420 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$1422 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1424 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1426 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1428 ;
  (* src = "sdram_controller.py:840" *)
  wire \$143 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1430 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1432 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1434 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1436 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1438 ;
  (* src = "sdram_controller.py:769" *)
  wire \$1440 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1442 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1444 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1446 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1448 ;
  (* src = "sdram_controller.py:849" *)
  wire \$145 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1450 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1452 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1454 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1456 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1458 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1460 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1462 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1464 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1466 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1468 ;
  (* src = "sdram_controller.py:869" *)
  wire \$147 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1470 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1472 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1474 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1476 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1478 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1480 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1482 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1484 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1486 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1488 ;
  (* src = "sdram_controller.py:915" *)
  wire \$149 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$1490 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1492 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1494 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1496 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1498 ;
  (* src = "sdram_controller.py:797" *)
  wire \$15 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1500 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1502 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1504 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1506 ;
  (* src = "sdram_controller.py:769" *)
  wire \$1508 ;
  (* src = "sdram_controller.py:917" *)
  wire \$151 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1510 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1512 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1514 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1516 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1518 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1520 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1522 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1524 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1526 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1528 ;
  (* src = "sdram_controller.py:926" *)
  wire \$153 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1530 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1532 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1534 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1536 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1538 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1540 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1542 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1544 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1546 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1548 ;
  (* src = "sdram_controller.py:955" *)
  wire \$155 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1550 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1552 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1554 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1556 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$1558 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1560 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1562 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1564 ;
  (* src = "sdram_controller.py:737" *)
  wire \$1566 ;
  (* src = "sdram_controller.py:374" *)
  wire \$1568 ;
  (* src = "sdram_controller.py:965" *)
  wire \$157 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1570 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1572 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1574 ;
  (* src = "sdram_controller.py:769" *)
  wire \$1576 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1578 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1580 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1582 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1584 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1586 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1588 ;
  (* src = "sdram_controller.py:970" *)
  wire \$159 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1590 ;
  (* src = "sdram_controller.py:917" *)
  wire \$1592 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1594 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1596 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1598 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1600 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1602 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1604 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1606 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1608 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$161 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1610 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$1612 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1614 ;
  (* src = "sdram_controller.py:355" *)
  wire \$1616 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1618 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1620 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1622 ;
  (* src = "sdram_controller.py:549" *)
  wire \$1624 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$1626 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1628 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$163 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1630 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1632 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1634 ;
  (* src = "sdram_controller.py:483" *)
  wire \$1636 ;
  (* src = "sdram_controller.py:754" *)
  wire \$1638 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1640 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1642 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1644 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1646 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1648 ;
  (* src = "sdram_controller.py:1020" *)
  wire \$165 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1650 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1652 ;
  (* src = "sdram_controller.py:837" *)
  wire \$1654 ;
  (* src = "sdram_controller.py:838" *)
  wire \$1656 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1658 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1660 ;
  (* src = "sdram_controller.py:440" *)
  wire \$1662 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1664 ;
  (* src = "sdram_controller.py:869" *)
  wire \$1666 ;
  (* src = "sdram_controller.py:915" *)
  wire \$1668 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$167 ;
  (* src = "sdram_controller.py:609" *)
  wire \$1670 ;
  (* src = "sdram_controller.py:610" *)
  wire \$1672 ;
  (* src = "sdram_controller.py:609" *)
  wire \$1674 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1676 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1678 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1680 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1682 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1684 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1686 ;
  (* src = "sdram_controller.py:970" *)
  wire \$1688 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$169 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$1690 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1692 ;
  (* src = "sdram_controller.py:396" *)
  wire \$1694 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1696 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$1698 ;
  (* src = "sdram_controller.py:795" *)
  wire \$17 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$1700 ;
  (* src = "sdram_controller.py:609" *)
  wire \$1702 ;
  (* src = "sdram_controller.py:610" *)
  wire \$1704 ;
  (* src = "sdram_controller.py:609" *)
  wire \$1706 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$1708 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$171 ;
  (* src = "sdram_controller.py:543" *)
  wire \$1710 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1712 ;
  (* src = "sdram_controller.py:748" *)
  wire \$1714 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1716 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1718 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1720 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1722 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1724 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1726 ;
  (* src = "sdram_controller.py:837" *)
  wire \$1728 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$173 ;
  (* src = "sdram_controller.py:838" *)
  wire \$1730 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1732 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1734 ;
  (* src = "sdram_controller.py:440" *)
  wire \$1736 ;
  (* src = "sdram_controller.py:439" *)
  wire \$1738 ;
  (* src = "sdram_controller.py:446" *)
  wire \$1740 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1742 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1744 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1746 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1748 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$175 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1750 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1752 ;
  (* src = "sdram_controller.py:970" *)
  wire \$1754 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$1756 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1758 ;
  (* src = "sdram_controller.py:396" *)
  wire \$1760 ;
  (* src = "sdram_controller.py:395" *)
  wire \$1762 ;
  (* src = "sdram_controller.py:402" *)
  wire \$1764 ;
  (* src = "sdram_controller.py:746" *)
  wire \$1766 ;
  (* src = "sdram_controller.py:769" *)
  wire \$1768 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$177 ;
  (* src = "sdram_controller.py:797" *)
  wire \$1770 ;
  (* src = "sdram_controller.py:932" *)
  wire \$1772 ;
  (* src = "sdram_controller.py:936" *)
  wire \$1774 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$1776 ;
  (* src = "sdram_controller.py:1082" *)
  wire \$1778 ;
  (* src = "sdram_controller.py:797" *)
  wire \$1780 ;
  (* src = "sdram_controller.py:814" *)
  wire \$1782 ;
  (* src = "sdram_controller.py:818" *)
  wire [9:0] \$1784 ;
  (* src = "sdram_controller.py:818" *)
  wire [10:0] \$1786 ;
  (* src = "sdram_controller.py:818" *)
  wire [11:0] \$1788 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$179 ;
  (* src = "sdram_controller.py:818" *)
  wire [12:0] \$1790 ;
  (* src = "sdram_controller.py:818" *)
  wire \$1792 ;
  (* src = "sdram_controller.py:951" *)
  wire \$1794 ;
  (* src = "sdram_controller.py:953" *)
  wire [9:0] \$1796 ;
  (* src = "sdram_controller.py:953" *)
  wire [10:0] \$1798 ;
  (* src = "sdram_controller.py:953" *)
  wire [11:0] \$1800 ;
  (* src = "sdram_controller.py:953" *)
  wire [12:0] \$1802 ;
  (* src = "sdram_controller.py:953" *)
  wire \$1804 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$1806 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1808 ;
  (* src = "sdram_controller.py:712" *)
  wire \$181 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1810 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1812 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1814 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1816 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1818 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1820 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1822 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1824 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1826 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1828 ;
  (* src = "sdram_controller.py:533" *)
  wire \$183 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1830 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1832 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1834 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1836 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1838 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1840 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1842 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1844 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1846 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1848 ;
  (* src = "sdram_controller.py:737" *)
  wire \$185 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1850 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1852 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1854 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1856 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1858 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1860 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1862 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1864 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1866 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1868 ;
  (* src = "sdram_controller.py:371" *)
  wire \$187 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1870 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1872 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1874 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1876 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1878 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1880 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1882 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1884 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1886 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1888 ;
  (* src = "sdram_controller.py:742" *)
  wire \$189 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1890 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1892 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1894 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1896 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1898 ;
  (* src = "sdram_controller.py:801" *)
  wire \$19 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1900 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1902 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1904 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1906 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1908 ;
  (* src = "sdram_controller.py:533" *)
  wire \$191 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1910 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1912 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1914 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1916 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1918 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1920 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1922 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1924 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1926 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1928 ;
  (* src = "sdram_controller.py:746" *)
  wire \$193 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1930 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1932 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1934 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1936 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1938 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1940 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1942 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1944 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1946 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1948 ;
  (* src = "sdram_controller.py:483" *)
  wire \$195 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1950 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1952 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1954 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1956 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1958 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1960 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1962 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1964 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1966 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1968 ;
  (* src = "sdram_controller.py:486" *)
  wire \$197 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1970 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1972 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1974 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1976 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1978 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1980 ;
  (* src = "sdram_controller.py:820" *)
  wire \$1982 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1984 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1986 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1988 ;
  (* src = "sdram_controller.py:754" *)
  wire \$199 ;
  (* src = "sdram_controller.py:327" *)
  wire \$1990 ;
  (* src = "sdram_controller.py:330" *)
  wire \$1992 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1994 ;
  (* src = "sdram_controller.py:955" *)
  wire \$1996 ;
  (* src = "sdram_controller.py:325" *)
  wire \$1998 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2000 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2002 ;
  (* src = "sdram_controller.py:327" *)
  wire \$2004 ;
  (* src = "sdram_controller.py:330" *)
  wire \$2006 ;
  (* src = "sdram_controller.py:334" *)
  wire \$2008 ;
  (* src = "sdram_controller.py:543" *)
  wire \$201 ;
  (* src = "sdram_controller.py:820" *)
  wire \$2010 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2012 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2014 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2016 ;
  (* src = "sdram_controller.py:327" *)
  wire \$2018 ;
  (* src = "sdram_controller.py:330" *)
  wire \$2020 ;
  (* src = "sdram_controller.py:334" *)
  wire \$2022 ;
  (* src = "sdram_controller.py:955" *)
  wire \$2024 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2026 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2028 ;
  (* src = "sdram_controller.py:546" *)
  wire \$203 ;
  (* src = "sdram_controller.py:325" *)
  wire \$2030 ;
  (* src = "sdram_controller.py:327" *)
  wire \$2032 ;
  (* src = "sdram_controller.py:330" *)
  wire \$2034 ;
  (* src = "sdram_controller.py:334" *)
  wire \$2036 ;
  (* src = "sdram_controller.py:820" *)
  wire \$2038 ;
  (* src = "sdram_controller.py:869" *)
  wire \$2040 ;
  (* src = "sdram_controller.py:915" *)
  wire \$2042 ;
  (* src = "sdram_controller.py:609" *)
  wire \$2044 ;
  (* src = "sdram_controller.py:610" *)
  wire \$2046 ;
  (* src = "sdram_controller.py:609" *)
  wire \$2048 ;
  (* src = "sdram_controller.py:549" *)
  wire \$205 ;
  (* src = "sdram_controller.py:616" *)
  wire \$2050 ;
  (* src = "sdram_controller.py:955" *)
  wire \$2052 ;
  (* src = "sdram_controller.py:970" *)
  wire \$2054 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$2056 ;
  (* src = "sdram_controller.py:395" *)
  wire \$2058 ;
  (* src = "sdram_controller.py:396" *)
  wire \$2060 ;
  (* src = "sdram_controller.py:395" *)
  wire \$2062 ;
  (* src = "sdram_controller.py:402" *)
  wire \$2064 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$2066 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$2068 ;
  (* src = "sdram_controller.py:758" *)
  wire \$207 ;
  (* src = "sdram_controller.py:609" *)
  wire \$2070 ;
  (* src = "sdram_controller.py:610" *)
  wire \$2072 ;
  (* src = "sdram_controller.py:609" *)
  wire \$2074 ;
  (* src = "sdram_controller.py:616" *)
  wire \$2076 ;
  (* src = "sdram_controller.py:837" *)
  wire \$2078 ;
  (* src = "sdram_controller.py:838" *)
  wire \$2080 ;
  (* src = "sdram_controller.py:840" *)
  wire \$2082 ;
  (* src = "sdram_controller.py:869" *)
  wire \$2084 ;
  (* src = "sdram_controller.py:910" *)
  wire \$2086 ;
  (* src = "sdram_controller.py:911" *)
  wire [8:0] \$2088 ;
  (* src = "sdram_controller.py:911" *)
  wire [8:0] \$2089 ;
  (* src = "sdram_controller.py:533" *)
  wire \$209 ;
  (* src = "sdram_controller.py:970" *)
  wire \$2091 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$2093 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$2095 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$2097 ;
  (* src = "sdram_controller.py:1053" *)
  wire [8:0] \$2099 ;
  (* src = "sdram_controller.py:820" *)
  wire \$21 ;
  (* src = "sdram_controller.py:1053" *)
  wire [8:0] \$2100 ;
  (* src = "sdram_controller.py:862" *)
  wire \$2102 ;
  (* src = "sdram_controller.py:917" *)
  wire \$2104 ;
  (* src = "sdram_controller.py:869" *)
  wire \$2106 ;
  (* src = "sdram_controller.py:917" *)
  wire \$2108 ;
  (* src = "sdram_controller.py:505" *)
  wire \$211 ;
  (* src = "sdram_controller.py:869" *)
  wire \$2110 ;
  (* src = "sdram_controller.py:917" *)
  wire \$2112 ;
  (* src = "sdram_controller.py:970" *)
  wire \$2114 ;
  (* src = "sdram_controller.py:997" *)
  wire \$2116 ;
  (* src = "sdram_controller.py:999" *)
  wire \$2118 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$2120 ;
  (* src = "sdram_controller.py:1061" *)
  wire \$2122 ;
  (* src = "sdram_controller.py:970" *)
  wire \$2124 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$2126 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$2128 ;
  (* src = "sdram_controller.py:820" *)
  wire \$213 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$2130 ;
  (* src = "sdram_controller.py:970" *)
  wire \$2132 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$2134 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$2136 ;
  (* src = "sdram_controller.py:970" *)
  wire \$2138 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$2140 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$2142 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$2144 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$2146 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$2148 ;
  (* src = "sdram_controller.py:325" *)
  wire \$215 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$2150 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$2152 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$2154 ;
  (* src = "sdram_controller.py:325" *)
  wire \$217 ;
  (* src = "sdram_controller.py:325" *)
  wire \$219 ;
  (* src = "sdram_controller.py:327" *)
  wire \$221 ;
  (* src = "sdram_controller.py:330" *)
  wire \$223 ;
  (* src = "sdram_controller.py:831" *)
  wire \$225 ;
  (* src = "sdram_controller.py:533" *)
  wire \$227 ;
  (* src = "sdram_controller.py:837" *)
  wire \$229 ;
  (* src = "sdram_controller.py:932" *)
  wire \$23 ;
  (* src = "sdram_controller.py:838" *)
  wire \$231 ;
  (* src = "sdram_controller.py:840" *)
  wire \$233 ;
  (* src = "sdram_controller.py:439" *)
  wire \$235 ;
  (* src = "sdram_controller.py:440" *)
  wire \$237 ;
  (* src = "sdram_controller.py:439" *)
  wire \$239 ;
  (* src = "sdram_controller.py:443" *)
  wire \$241 ;
  (* src = "sdram_controller.py:849" *)
  wire \$243 ;
  (* src = "sdram_controller.py:533" *)
  wire \$245 ;
  (* src = "sdram_controller.py:869" *)
  wire \$247 ;
  (* src = "sdram_controller.py:915" *)
  wire \$249 ;
  (* src = "sdram_controller.py:936" *)
  wire \$25 ;
  (* src = "sdram_controller.py:609" *)
  wire \$251 ;
  (* src = "sdram_controller.py:610" *)
  wire \$253 ;
  (* src = "sdram_controller.py:609" *)
  wire \$255 ;
  (* src = "sdram_controller.py:613" *)
  wire \$257 ;
  (* src = "sdram_controller.py:917" *)
  wire \$259 ;
  (* src = "sdram_controller.py:352" *)
  wire \$261 ;
  (* src = "sdram_controller.py:926" *)
  wire \$263 ;
  (* src = "sdram_controller.py:533" *)
  wire \$265 ;
  (* src = "sdram_controller.py:955" *)
  wire \$267 ;
  (* src = "sdram_controller.py:325" *)
  wire \$269 ;
  (* src = "sdram_controller.py:955" *)
  wire \$27 ;
  (* src = "sdram_controller.py:325" *)
  wire \$271 ;
  (* src = "sdram_controller.py:325" *)
  wire \$273 ;
  (* src = "sdram_controller.py:327" *)
  wire \$275 ;
  (* src = "sdram_controller.py:330" *)
  wire \$277 ;
  (* src = "sdram_controller.py:965" *)
  wire \$279 ;
  (* src = "sdram_controller.py:505" *)
  wire \$281 ;
  (* src = "sdram_controller.py:970" *)
  wire \$283 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$285 ;
  (* src = "sdram_controller.py:395" *)
  wire \$287 ;
  (* src = "sdram_controller.py:396" *)
  wire \$289 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$29 ;
  (* src = "sdram_controller.py:395" *)
  wire \$291 ;
  (* src = "sdram_controller.py:399" *)
  wire \$293 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$295 ;
  (* src = "sdram_controller.py:1020" *)
  wire \$297 ;
  (* src = "sdram_controller.py:533" *)
  wire \$299 ;
  (* src = "sdram_controller.py:655" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$301 ;
  (* src = "sdram_controller.py:609" *)
  wire \$303 ;
  (* src = "sdram_controller.py:610" *)
  wire \$305 ;
  (* src = "sdram_controller.py:609" *)
  wire \$307 ;
  (* src = "sdram_controller.py:613" *)
  wire \$309 ;
  (* src = "sdram_controller.py:1082" *)
  wire \$31 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$311 ;
  (* src = "sdram_controller.py:533" *)
  wire \$313 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$315 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$317 ;
  (* src = "sdram_controller.py:352" *)
  wire \$319 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$321 ;
  (* src = "sdram_controller.py:533" *)
  wire \$323 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$325 ;
  (* src = "sdram_controller.py:543" *)
  wire \$327 ;
  (* src = "sdram_controller.py:546" *)
  wire \$329 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$33 ;
  (* src = "sdram_controller.py:549" *)
  wire \$331 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$333 ;
  (* src = "sdram_controller.py:533" *)
  wire \$335 ;
  (* src = "sdram_controller.py:712" *)
  wire \$337 ;
  (* src = "sdram_controller.py:533" *)
  wire \$339 ;
  (* src = "sdram_controller.py:536" *)
  wire \$341 ;
  (* src = "sdram_controller.py:737" *)
  wire \$343 ;
  (* src = "sdram_controller.py:371" *)
  wire \$345 ;
  (* src = "sdram_controller.py:374" *)
  wire \$347 ;
  (* src = "sdram_controller.py:742" *)
  wire \$349 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$35 ;
  (* src = "sdram_controller.py:533" *)
  wire \$351 ;
  (* src = "sdram_controller.py:536" *)
  wire \$353 ;
  (* src = "sdram_controller.py:746" *)
  wire \$355 ;
  (* src = "sdram_controller.py:483" *)
  wire \$357 ;
  (* src = "sdram_controller.py:486" *)
  wire \$359 ;
  (* src = "sdram_controller.py:489" *)
  wire \$361 ;
  (* src = "sdram_controller.py:754" *)
  wire \$363 ;
  (* src = "sdram_controller.py:543" *)
  wire \$365 ;
  (* src = "sdram_controller.py:546" *)
  wire \$367 ;
  (* src = "sdram_controller.py:549" *)
  wire \$369 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$37 ;
  (* src = "sdram_controller.py:758" *)
  wire \$371 ;
  (* src = "sdram_controller.py:533" *)
  wire \$373 ;
  (* src = "sdram_controller.py:536" *)
  wire \$375 ;
  (* src = "sdram_controller.py:505" *)
  wire \$377 ;
  (* src = "sdram_controller.py:508" *)
  wire \$379 ;
  (* src = "sdram_controller.py:820" *)
  wire \$381 ;
  (* src = "sdram_controller.py:325" *)
  wire \$383 ;
  (* src = "sdram_controller.py:325" *)
  wire \$385 ;
  (* src = "sdram_controller.py:325" *)
  wire \$387 ;
  (* src = "sdram_controller.py:327" *)
  wire \$389 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$39 ;
  (* src = "sdram_controller.py:330" *)
  wire \$391 ;
  (* src = "sdram_controller.py:831" *)
  wire \$393 ;
  (* src = "sdram_controller.py:533" *)
  wire \$395 ;
  (* src = "sdram_controller.py:536" *)
  wire \$397 ;
  (* src = "sdram_controller.py:837" *)
  wire \$399 ;
  (* src = "sdram_controller.py:838" *)
  wire \$401 ;
  (* src = "sdram_controller.py:840" *)
  wire \$403 ;
  (* src = "sdram_controller.py:439" *)
  wire \$405 ;
  (* src = "sdram_controller.py:440" *)
  wire \$407 ;
  (* src = "sdram_controller.py:439" *)
  wire \$409 ;
  (* src = "sdram_controller.py:1110" *)
  wire \$41 ;
  (* src = "sdram_controller.py:443" *)
  wire \$411 ;
  (* src = "sdram_controller.py:446" *)
  wire \$413 ;
  (* src = "sdram_controller.py:849" *)
  wire \$415 ;
  (* src = "sdram_controller.py:533" *)
  wire \$417 ;
  (* src = "sdram_controller.py:536" *)
  wire \$419 ;
  (* src = "sdram_controller.py:869" *)
  wire \$421 ;
  (* src = "sdram_controller.py:915" *)
  wire \$423 ;
  (* src = "sdram_controller.py:609" *)
  wire \$425 ;
  (* src = "sdram_controller.py:610" *)
  wire \$427 ;
  (* src = "sdram_controller.py:609" *)
  wire \$429 ;
  (* src = "sdram_controller.py:1112" *)
  wire \$43 ;
  (* src = "sdram_controller.py:613" *)
  wire \$431 ;
  (* src = "sdram_controller.py:616" *)
  wire \$433 ;
  (* src = "sdram_controller.py:917" *)
  wire \$435 ;
  (* src = "sdram_controller.py:352" *)
  wire \$437 ;
  (* src = "sdram_controller.py:355" *)
  wire \$439 ;
  (* src = "sdram_controller.py:926" *)
  wire \$441 ;
  (* src = "sdram_controller.py:533" *)
  wire \$443 ;
  (* src = "sdram_controller.py:536" *)
  wire \$445 ;
  (* src = "sdram_controller.py:955" *)
  wire \$447 ;
  (* src = "sdram_controller.py:325" *)
  wire \$449 ;
  (* src = "sdram_controller.py:722" *)
  wire \$45 ;
  (* src = "sdram_controller.py:325" *)
  wire \$451 ;
  (* src = "sdram_controller.py:325" *)
  wire \$453 ;
  (* src = "sdram_controller.py:327" *)
  wire \$455 ;
  (* src = "sdram_controller.py:330" *)
  wire \$457 ;
  (* src = "sdram_controller.py:965" *)
  wire \$459 ;
  (* src = "sdram_controller.py:505" *)
  wire \$461 ;
  (* src = "sdram_controller.py:508" *)
  wire \$463 ;
  (* src = "sdram_controller.py:970" *)
  wire \$465 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$467 ;
  (* src = "sdram_controller.py:395" *)
  wire \$469 ;
  (* src = "sdram_controller.py:723" *)
  wire \$47 ;
  (* src = "sdram_controller.py:396" *)
  wire \$471 ;
  (* src = "sdram_controller.py:395" *)
  wire \$473 ;
  (* src = "sdram_controller.py:399" *)
  wire \$475 ;
  (* src = "sdram_controller.py:402" *)
  wire \$477 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$479 ;
  (* src = "sdram_controller.py:1020" *)
  wire \$481 ;
  (* src = "sdram_controller.py:533" *)
  wire \$483 ;
  (* src = "sdram_controller.py:536" *)
  wire \$485 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$487 ;
  (* src = "sdram_controller.py:609" *)
  wire \$489 ;
  (* src = "sdram_controller.py:769" *)
  wire \$49 ;
  (* src = "sdram_controller.py:610" *)
  wire \$491 ;
  (* src = "sdram_controller.py:609" *)
  wire \$493 ;
  (* src = "sdram_controller.py:613" *)
  wire \$495 ;
  (* src = "sdram_controller.py:616" *)
  wire \$497 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$499 ;
  (* src = "sdram_controller.py:655" *)
  wire \$5 ;
  (* src = "sdram_controller.py:533" *)
  wire \$501 ;
  (* src = "sdram_controller.py:536" *)
  wire \$503 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$505 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$507 ;
  (* src = "sdram_controller.py:352" *)
  wire \$509 ;
  (* src = "sdram_controller.py:797" *)
  wire \$51 ;
  (* src = "sdram_controller.py:355" *)
  wire \$511 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$513 ;
  (* src = "sdram_controller.py:533" *)
  wire \$515 ;
  (* src = "sdram_controller.py:536" *)
  wire \$517 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$519 ;
  (* src = "sdram_controller.py:543" *)
  wire \$521 ;
  (* src = "sdram_controller.py:546" *)
  wire \$523 ;
  (* src = "sdram_controller.py:549" *)
  wire \$525 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$527 ;
  (* src = "sdram_controller.py:533" *)
  wire \$529 ;
  (* src = "sdram_controller.py:820" *)
  wire \$53 ;
  (* src = "sdram_controller.py:536" *)
  wire \$531 ;
  (* src = "sdram_controller.py:712" *)
  wire \$533 ;
  (* src = "sdram_controller.py:536" *)
  wire \$535 ;
  (* src = "sdram_controller.py:737" *)
  wire \$537 ;
  (* src = "sdram_controller.py:386" *)
  wire \$539 ;
  (* src = "sdram_controller.py:388" *)
  wire \$541 ;
  (* src = "sdram_controller.py:742" *)
  wire \$543 ;
  (* src = "sdram_controller.py:536" *)
  wire \$545 ;
  (* src = "sdram_controller.py:746" *)
  wire \$547 ;
  (* src = "sdram_controller.py:483" *)
  wire \$549 ;
  (* src = "sdram_controller.py:955" *)
  wire \$55 ;
  (* src = "sdram_controller.py:497" *)
  wire \$551 ;
  (* src = "sdram_controller.py:499" *)
  wire \$553 ;
  (* src = "sdram_controller.py:754" *)
  wire \$555 ;
  (* src = "sdram_controller.py:543" *)
  wire \$557 ;
  (* src = "sdram_controller.py:549" *)
  wire \$559 ;
  (* src = "sdram_controller.py:758" *)
  wire \$561 ;
  (* src = "sdram_controller.py:536" *)
  wire \$563 ;
  (* src = "sdram_controller.py:508" *)
  wire \$565 ;
  (* src = "sdram_controller.py:820" *)
  wire \$567 ;
  (* src = "sdram_controller.py:325" *)
  wire \$569 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$57 ;
  (* src = "sdram_controller.py:325" *)
  wire \$571 ;
  (* src = "sdram_controller.py:325" *)
  wire \$573 ;
  (* src = "sdram_controller.py:327" *)
  wire \$575 ;
  (* src = "sdram_controller.py:330" *)
  wire \$577 ;
  (* src = "sdram_controller.py:831" *)
  wire \$579 ;
  (* src = "sdram_controller.py:536" *)
  wire \$581 ;
  (* src = "sdram_controller.py:837" *)
  wire \$583 ;
  (* src = "sdram_controller.py:838" *)
  wire \$585 ;
  (* src = "sdram_controller.py:840" *)
  wire \$587 ;
  (* src = "sdram_controller.py:439" *)
  wire \$589 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$59 ;
  (* src = "sdram_controller.py:440" *)
  wire \$591 ;
  (* src = "sdram_controller.py:439" *)
  wire \$593 ;
  (* src = "sdram_controller.py:446" *)
  wire \$595 ;
  (* src = "sdram_controller.py:849" *)
  wire \$597 ;
  (* src = "sdram_controller.py:536" *)
  wire \$599 ;
  (* src = "sdram_controller.py:869" *)
  wire \$601 ;
  (* src = "sdram_controller.py:915" *)
  wire \$603 ;
  (* src = "sdram_controller.py:609" *)
  wire \$605 ;
  (* src = "sdram_controller.py:610" *)
  wire \$607 ;
  (* src = "sdram_controller.py:609" *)
  wire \$609 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$61 ;
  (* src = "sdram_controller.py:616" *)
  wire \$611 ;
  (* src = "sdram_controller.py:917" *)
  wire \$613 ;
  (* src = "sdram_controller.py:355" *)
  wire \$615 ;
  (* src = "sdram_controller.py:926" *)
  wire \$617 ;
  (* src = "sdram_controller.py:536" *)
  wire \$619 ;
  (* src = "sdram_controller.py:955" *)
  wire \$621 ;
  (* src = "sdram_controller.py:325" *)
  wire \$623 ;
  (* src = "sdram_controller.py:325" *)
  wire \$625 ;
  (* src = "sdram_controller.py:325" *)
  wire \$627 ;
  (* src = "sdram_controller.py:327" *)
  wire \$629 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$63 ;
  (* src = "sdram_controller.py:330" *)
  wire \$631 ;
  (* src = "sdram_controller.py:965" *)
  wire \$633 ;
  (* src = "sdram_controller.py:508" *)
  wire \$635 ;
  (* src = "sdram_controller.py:970" *)
  wire \$637 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$639 ;
  (* src = "sdram_controller.py:395" *)
  wire \$641 ;
  (* src = "sdram_controller.py:396" *)
  wire \$643 ;
  (* src = "sdram_controller.py:395" *)
  wire \$645 ;
  (* src = "sdram_controller.py:402" *)
  wire \$647 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$649 ;
  (* src = "sdram_controller.py:712" *)
  wire \$65 ;
  (* src = "sdram_controller.py:1020" *)
  wire \$651 ;
  (* src = "sdram_controller.py:536" *)
  wire \$653 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$655 ;
  (* src = "sdram_controller.py:609" *)
  wire \$657 ;
  (* src = "sdram_controller.py:610" *)
  wire \$659 ;
  (* src = "sdram_controller.py:609" *)
  wire \$661 ;
  (* src = "sdram_controller.py:616" *)
  wire \$663 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$665 ;
  (* src = "sdram_controller.py:536" *)
  wire \$667 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$669 ;
  (* src = "sdram_controller.py:737" *)
  wire \$67 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$671 ;
  (* src = "sdram_controller.py:355" *)
  wire \$673 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$675 ;
  (* src = "sdram_controller.py:536" *)
  wire \$677 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$679 ;
  (* src = "sdram_controller.py:543" *)
  wire \$681 ;
  (* src = "sdram_controller.py:549" *)
  wire \$683 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$685 ;
  (* src = "sdram_controller.py:536" *)
  wire \$687 ;
  (* src = "sdram_controller.py:712" *)
  wire \$689 ;
  (* src = "sdram_controller.py:742" *)
  wire \$69 ;
  (* src = "sdram_controller.py:536" *)
  wire \$691 ;
  (* src = "sdram_controller.py:737" *)
  wire \$693 ;
  (* src = "sdram_controller.py:374" *)
  wire \$695 ;
  (* src = "sdram_controller.py:742" *)
  wire \$697 ;
  (* src = "sdram_controller.py:536" *)
  wire \$699 ;
  (* src = "sdram_controller.py:655" *)
  wire \$7 ;
  (* src = "sdram_controller.py:746" *)
  wire \$701 ;
  (* src = "sdram_controller.py:483" *)
  wire \$703 ;
  (* src = "sdram_controller.py:489" *)
  wire \$705 ;
  (* src = "sdram_controller.py:754" *)
  wire \$707 ;
  (* src = "sdram_controller.py:543" *)
  wire \$709 ;
  (* src = "sdram_controller.py:746" *)
  wire \$71 ;
  (* src = "sdram_controller.py:549" *)
  wire \$711 ;
  (* src = "sdram_controller.py:758" *)
  wire \$713 ;
  (* src = "sdram_controller.py:536" *)
  wire \$715 ;
  (* src = "sdram_controller.py:508" *)
  wire \$717 ;
  (* src = "sdram_controller.py:820" *)
  wire \$719 ;
  (* src = "sdram_controller.py:325" *)
  wire \$721 ;
  (* src = "sdram_controller.py:325" *)
  wire \$723 ;
  (* src = "sdram_controller.py:325" *)
  wire \$725 ;
  (* src = "sdram_controller.py:327" *)
  wire \$727 ;
  (* src = "sdram_controller.py:330" *)
  wire \$729 ;
  (* src = "sdram_controller.py:754" *)
  wire \$73 ;
  (* src = "sdram_controller.py:831" *)
  wire \$731 ;
  (* src = "sdram_controller.py:536" *)
  wire \$733 ;
  (* src = "sdram_controller.py:837" *)
  wire \$735 ;
  (* src = "sdram_controller.py:838" *)
  wire \$737 ;
  (* src = "sdram_controller.py:840" *)
  wire \$739 ;
  (* src = "sdram_controller.py:439" *)
  wire \$741 ;
  (* src = "sdram_controller.py:440" *)
  wire \$743 ;
  (* src = "sdram_controller.py:439" *)
  wire \$745 ;
  (* src = "sdram_controller.py:446" *)
  wire \$747 ;
  (* src = "sdram_controller.py:849" *)
  wire \$749 ;
  (* src = "sdram_controller.py:758" *)
  wire \$75 ;
  (* src = "sdram_controller.py:536" *)
  wire \$751 ;
  (* src = "sdram_controller.py:917" *)
  wire \$753 ;
  (* src = "sdram_controller.py:355" *)
  wire \$755 ;
  (* src = "sdram_controller.py:926" *)
  wire \$757 ;
  (* src = "sdram_controller.py:536" *)
  wire \$759 ;
  (* src = "sdram_controller.py:955" *)
  wire \$761 ;
  (* src = "sdram_controller.py:325" *)
  wire \$763 ;
  (* src = "sdram_controller.py:325" *)
  wire \$765 ;
  (* src = "sdram_controller.py:325" *)
  wire \$767 ;
  (* src = "sdram_controller.py:327" *)
  wire \$769 ;
  (* src = "sdram_controller.py:820" *)
  wire \$77 ;
  (* src = "sdram_controller.py:330" *)
  wire \$771 ;
  (* src = "sdram_controller.py:965" *)
  wire \$773 ;
  (* src = "sdram_controller.py:508" *)
  wire \$775 ;
  (* src = "sdram_controller.py:970" *)
  wire \$777 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$779 ;
  (* src = "sdram_controller.py:395" *)
  wire \$781 ;
  (* src = "sdram_controller.py:396" *)
  wire \$783 ;
  (* src = "sdram_controller.py:395" *)
  wire \$785 ;
  (* src = "sdram_controller.py:402" *)
  wire \$787 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$789 ;
  (* src = "sdram_controller.py:831" *)
  wire \$79 ;
  (* src = "sdram_controller.py:1020" *)
  wire \$791 ;
  (* src = "sdram_controller.py:536" *)
  wire \$793 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$795 ;
  (* src = "sdram_controller.py:536" *)
  wire \$797 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$799 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$801 ;
  (* src = "sdram_controller.py:355" *)
  wire \$803 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$805 ;
  (* src = "sdram_controller.py:536" *)
  wire \$807 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$809 ;
  (* src = "sdram_controller.py:837" *)
  wire \$81 ;
  (* src = "sdram_controller.py:543" *)
  wire \$811 ;
  (* src = "sdram_controller.py:549" *)
  wire \$813 ;
  (* src = "sdram_controller.py:1099" *)
  wire \$815 ;
  (* src = "sdram_controller.py:536" *)
  wire \$817 ;
  (* src = "sdram_controller.py:712" *)
  wire \$819 ;
  (* src = "sdram_controller.py:737" *)
  wire \$821 ;
  (* src = "sdram_controller.py:769" *)
  wire \$823 ;
  (* src = "sdram_controller.py:712" *)
  wire \$825 ;
  (* src = "sdram_controller.py:722" *)
  wire \$827 ;
  (* src = "sdram_controller.py:723" *)
  wire \$829 ;
  (* src = "sdram_controller.py:838" *)
  wire \$83 ;
  (* src = "sdram_controller.py:724" *)
  wire [15:0] \$831 ;
  (* src = "sdram_controller.py:724" *)
  wire [15:0] \$832 ;
  (* src = "sdram_controller.py:712" *)
  wire \$834 ;
  (* src = "sdram_controller.py:722" *)
  wire \$836 ;
  (* src = "sdram_controller.py:723" *)
  wire \$838 ;
  (* src = "sdram_controller.py:737" *)
  wire \$840 ;
  (* src = "sdram_controller.py:742" *)
  wire \$842 ;
  (* src = "sdram_controller.py:746" *)
  wire \$844 ;
  (* src = "sdram_controller.py:754" *)
  wire \$846 ;
  (* src = "sdram_controller.py:758" *)
  wire \$848 ;
  (* src = "sdram_controller.py:840" *)
  wire \$85 ;
  (* src = "sdram_controller.py:763" *)
  wire \$850 ;
  (* src = "sdram_controller.py:764" *)
  wire \$852 ;
  (* src = "sdram_controller.py:766" *)
  wire \$854 ;
  (* src = "sdram_controller.py:769" *)
  wire \$856 ;
  (* src = "sdram_controller.py:814" *)
  wire \$858 ;
  (* src = "sdram_controller.py:820" *)
  wire \$860 ;
  (* src = "sdram_controller.py:831" *)
  wire \$862 ;
  (* src = "sdram_controller.py:837" *)
  wire \$864 ;
  (* src = "sdram_controller.py:838" *)
  wire \$866 ;
  (* src = "sdram_controller.py:840" *)
  wire \$868 ;
  (* src = "sdram_controller.py:849" *)
  wire \$87 ;
  (* src = "sdram_controller.py:849" *)
  wire \$870 ;
  (* src = "sdram_controller.py:853" *)
  wire \$872 ;
  (* src = "sdram_controller.py:862" *)
  wire \$874 ;
  (* src = "sdram_controller.py:869" *)
  wire \$876 ;
  (* src = "sdram_controller.py:910" *)
  wire \$878 ;
  (* src = "sdram_controller.py:917" *)
  wire \$880 ;
  (* src = "sdram_controller.py:926" *)
  wire \$882 ;
  (* src = "sdram_controller.py:932" *)
  wire \$884 ;
  (* src = "sdram_controller.py:936" *)
  wire \$886 ;
  (* src = "sdram_controller.py:951" *)
  wire \$888 ;
  (* src = "sdram_controller.py:869" *)
  wire \$89 ;
  (* src = "sdram_controller.py:955" *)
  wire \$890 ;
  (* src = "sdram_controller.py:965" *)
  wire \$892 ;
  (* src = "sdram_controller.py:970" *)
  wire \$894 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$896 ;
  (* src = "sdram_controller.py:1013" *)
  wire \$898 ;
  (* src = "sdram_controller.py:722" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1052" *)
  wire \$900 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$902 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$904 ;
  (* src = "sdram_controller.py:1078" *)
  wire \$906 ;
  (* src = "sdram_controller.py:1082" *)
  wire \$908 ;
  (* src = "sdram_controller.py:915" *)
  wire \$91 ;
  (* src = "sdram_controller.py:712" *)
  wire \$910 ;
  (* src = "sdram_controller.py:737" *)
  wire \$912 ;
  (* src = "sdram_controller.py:374" *)
  wire \$914 ;
  (* src = "sdram_controller.py:746" *)
  wire \$916 ;
  (* src = "sdram_controller.py:483" *)
  wire \$918 ;
  (* src = "sdram_controller.py:489" *)
  wire \$920 ;
  (* src = "sdram_controller.py:754" *)
  wire \$922 ;
  (* src = "sdram_controller.py:543" *)
  wire \$924 ;
  (* src = "sdram_controller.py:549" *)
  wire \$926 ;
  (* src = "sdram_controller.py:508" *)
  wire \$928 ;
  (* src = "sdram_controller.py:917" *)
  wire \$93 ;
  (* src = "sdram_controller.py:820" *)
  wire \$930 ;
  (* src = "sdram_controller.py:325" *)
  wire \$932 ;
  (* src = "sdram_controller.py:325" *)
  wire \$934 ;
  (* src = "sdram_controller.py:325" *)
  wire \$936 ;
  (* src = "sdram_controller.py:327" *)
  wire \$938 ;
  (* src = "sdram_controller.py:330" *)
  wire \$940 ;
  (* src = "sdram_controller.py:837" *)
  wire \$942 ;
  (* src = "sdram_controller.py:838" *)
  wire \$944 ;
  (* src = "sdram_controller.py:840" *)
  wire \$946 ;
  (* src = "sdram_controller.py:439" *)
  wire \$948 ;
  (* src = "sdram_controller.py:926" *)
  wire \$95 ;
  (* src = "sdram_controller.py:440" *)
  wire \$950 ;
  (* src = "sdram_controller.py:439" *)
  wire \$952 ;
  (* src = "sdram_controller.py:446" *)
  wire \$954 ;
  (* src = "sdram_controller.py:917" *)
  wire \$956 ;
  (* src = "sdram_controller.py:355" *)
  wire \$958 ;
  (* src = "sdram_controller.py:955" *)
  wire \$960 ;
  (* src = "sdram_controller.py:325" *)
  wire \$962 ;
  (* src = "sdram_controller.py:325" *)
  wire \$964 ;
  (* src = "sdram_controller.py:325" *)
  wire \$966 ;
  (* src = "sdram_controller.py:327" *)
  wire \$968 ;
  (* src = "sdram_controller.py:955" *)
  wire \$97 ;
  (* src = "sdram_controller.py:330" *)
  wire \$970 ;
  (* src = "sdram_controller.py:965" *)
  wire \$972 ;
  (* src = "sdram_controller.py:508" *)
  wire \$974 ;
  (* src = "sdram_controller.py:970" *)
  wire \$976 ;
  (* src = "sdram_controller.py:1001" *)
  wire \$978 ;
  (* src = "sdram_controller.py:395" *)
  wire \$980 ;
  (* src = "sdram_controller.py:396" *)
  wire \$982 ;
  (* src = "sdram_controller.py:395" *)
  wire \$984 ;
  (* src = "sdram_controller.py:402" *)
  wire \$986 ;
  (* src = "sdram_controller.py:1069" *)
  wire \$988 ;
  (* src = "sdram_controller.py:965" *)
  wire \$99 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$990 ;
  (* src = "sdram_controller.py:355" *)
  wire \$992 ;
  (* src = "sdram_controller.py:1094" *)
  wire \$994 ;
  (* src = "sdram_controller.py:543" *)
  wire \$996 ;
  (* src = "sdram_controller.py:549" *)
  wire \$998 ;
  (* src = "sdram_controller.py:235" *)
  reg allBanksIdle;
  (* src = "sdram_controller.py:1177" *)
  reg bankController0_bankActivated;
  (* src = "sdram_controller.py:1176" *)
  wire bankController0_bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  wire bankController0_bankCanPreCharge;
  (* src = "sdram_controller.py:1169" *)
  wire [9:0] bankController0_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1174" *)
  wire bankController0_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankController0_bankState = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankController0_bankState$next ;
  (* src = "sdram_controller.py:1178" *)
  reg bankController0_otherBankActivated;
  (* src = "sdram_controller.py:1177" *)
  reg bankController1_bankActivated;
  (* src = "sdram_controller.py:1176" *)
  wire bankController1_bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  wire bankController1_bankCanPreCharge;
  (* src = "sdram_controller.py:1169" *)
  wire [9:0] bankController1_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1174" *)
  wire bankController1_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankController1_bankState = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankController1_bankState$next ;
  (* src = "sdram_controller.py:1178" *)
  reg bankController1_otherBankActivated;
  (* src = "sdram_controller.py:1177" *)
  reg bankController2_bankActivated;
  (* src = "sdram_controller.py:1176" *)
  wire bankController2_bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  wire bankController2_bankCanPreCharge;
  (* src = "sdram_controller.py:1169" *)
  wire [9:0] bankController2_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1174" *)
  wire bankController2_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankController2_bankState = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankController2_bankState$next ;
  (* src = "sdram_controller.py:1178" *)
  reg bankController2_otherBankActivated;
  (* src = "sdram_controller.py:1177" *)
  reg bankController3_bankActivated;
  (* src = "sdram_controller.py:1176" *)
  wire bankController3_bankCanActivate;
  (* src = "sdram_controller.py:1175" *)
  wire bankController3_bankCanPreCharge;
  (* src = "sdram_controller.py:1169" *)
  wire [9:0] bankController3_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1174" *)
  wire bankController3_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankController3_bankState = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankController3_bankState$next ;
  (* src = "sdram_controller.py:1178" *)
  reg bankController3_otherBankActivated;
  (* src = "sdram_controller.py:234" *)
  reg banksShouldRefresh;
  (* src = "sdram_controller.py:257" *)
  reg burstWritesMode = 1'h0;
  (* src = "sdram_controller.py:257" *)
  reg \burstWritesMode$next ;
  (* src = "sdram_controller.py:1288" *)
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1288" *)
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:250" *)
  reg cmdCompleted;
  (* src = "sdram_controller.py:251" *)
  reg [3:0] cmdIndex = 4'h0;
  (* src = "sdram_controller.py:251" *)
  reg [3:0] \cmdIndex$next ;
  (* src = "sdram_controller.py:249" *)
  reg [1:0] cmdRemainingCyclesCounter;
  (* src = "sdram_controller.py:245" *)
  reg [20:0] ctrlAddress = 21'h000000;
  (* src = "sdram_controller.py:245" *)
  reg [20:0] \ctrlAddress$next ;
  (* src = "sdram_controller.py:218" *)
  input ctrlRd;
  wire ctrlRd;
  (* src = "sdram_controller.py:217" *)
  input [20:0] ctrlRdAddress;
  wire [20:0] ctrlRdAddress;
  (* src = "sdram_controller.py:219" *)
  output [23:0] ctrlRdDataOut;
  reg [23:0] ctrlRdDataOut;
  (* src = "sdram_controller.py:221" *)
  reg ctrlRdInProgress = 1'h0;
  (* src = "sdram_controller.py:221" *)
  reg \ctrlRdInProgress$next ;
  (* src = "sdram_controller.py:220" *)
  output ctrlRdIncAddress;
  reg ctrlRdIncAddress = 1'h0;
  (* src = "sdram_controller.py:220" *)
  reg \ctrlRdIncAddress$next ;
  (* src = "sdram_controller.py:209" *)
  output ctrlReady;
  reg ctrlReady = 1'h0;
  (* src = "sdram_controller.py:209" *)
  reg \ctrlReady$next ;
  (* src = "sdram_controller.py:212" *)
  input ctrlWr;
  wire ctrlWr;
  (* src = "sdram_controller.py:211" *)
  input [20:0] ctrlWrAddress;
  wire [20:0] ctrlWrAddress;
  (* src = "sdram_controller.py:213" *)
  input [23:0] ctrlWrDataIn;
  wire [23:0] ctrlWrDataIn;
  (* src = "sdram_controller.py:215" *)
  reg ctrlWrInProgress = 1'h0;
  (* src = "sdram_controller.py:215" *)
  reg \ctrlWrInProgress$next ;
  (* src = "sdram_controller.py:214" *)
  output ctrlWrIncAddress;
  reg ctrlWrIncAddress = 1'h0;
  (* src = "sdram_controller.py:214" *)
  reg \ctrlWrIncAddress$next ;
  (* enum_base_type = "Command" *)
  (* enum_value_00000 = "NoCommand" *)
  (* enum_value_00001 = "BankActivate" *)
  (* enum_value_00010 = "BankPreCharge" *)
  (* enum_value_00011 = "PreChargeAll" *)
  (* enum_value_00100 = "Write" *)
  (* enum_value_00101 = "WriteAndAutoPreCharge" *)
  (* enum_value_00110 = "Read" *)
  (* enum_value_00111 = "ReadAndAutoPreCharge" *)
  (* enum_value_01000 = "ModeRegisterSet" *)
  (* enum_value_01001 = "NoOperation" *)
  (* enum_value_01010 = "BurstStop" *)
  (* enum_value_01011 = "DeviceDeSelect" *)
  (* enum_value_01100 = "AutoRefresh" *)
  (* enum_value_01101 = "SelfRefreshEntry" *)
  (* enum_value_01110 = "SelfRefreshExit" *)
  (* enum_value_01111 = "ClockSuspendModeExit" *)
  (* enum_value_10000 = "PowerDownModeExit" *)
  (* enum_value_10001 = "DataWrite_OutputEnable" *)
  (* enum_value_10010 = "DataMask_OutputDisable" *)
  (* src = "sdram_controller.py:248" *)
  reg [4:0] currentCommand = 5'h00;
  (* src = "sdram_controller.py:248" *)
  reg [4:0] \currentCommand$next ;
  (* enum_base_type = "SDRAMControllerStates" *)
  (* enum_value_000 = "InitOp" *)
  (* enum_value_001 = "ConfigurationOp" *)
  (* enum_value_010 = "Idle" *)
  (* enum_value_011 = "RefreshOp" *)
  (* enum_value_100 = "WriteBurstOp" *)
  (* enum_value_101 = "WriteOp" *)
  (* enum_value_110 = "ReadOp" *)
  (* enum_value_111 = "Error" *)
  (* src = "sdram_controller.py:226" *)
  reg [2:0] currentControllerState;
  (* src = "sdram_controller.py:255" *)
  reg [3:0] delayCounter = 4'h0;
  (* src = "sdram_controller.py:255" *)
  reg [3:0] \delayCounter$next ;
  (* src = "sdram_controller.py:224" *)
  reg errorState = 1'h0;
  (* src = "sdram_controller.py:224" *)
  reg \errorState$next ;
  (* enum_base_type = "Command" *)
  (* enum_value_00000 = "NoCommand" *)
  (* enum_value_00001 = "BankActivate" *)
  (* enum_value_00010 = "BankPreCharge" *)
  (* enum_value_00011 = "PreChargeAll" *)
  (* enum_value_00100 = "Write" *)
  (* enum_value_00101 = "WriteAndAutoPreCharge" *)
  (* enum_value_00110 = "Read" *)
  (* enum_value_00111 = "ReadAndAutoPreCharge" *)
  (* enum_value_01000 = "ModeRegisterSet" *)
  (* enum_value_01001 = "NoOperation" *)
  (* enum_value_01010 = "BurstStop" *)
  (* enum_value_01011 = "DeviceDeSelect" *)
  (* enum_value_01100 = "AutoRefresh" *)
  (* enum_value_01101 = "SelfRefreshEntry" *)
  (* enum_value_01110 = "SelfRefreshExit" *)
  (* enum_value_01111 = "ClockSuspendModeExit" *)
  (* enum_value_10000 = "PowerDownModeExit" *)
  (* enum_value_10001 = "DataWrite_OutputEnable" *)
  (* enum_value_10010 = "DataMask_OutputDisable" *)
  (* src = "sdram_controller.py:247" *)
  reg [4:0] nextCommand;
  (* src = "sdram_controller.py:258" *)
  reg [7:0] pageColumnIndex = 8'h00;
  (* src = "sdram_controller.py:258" *)
  reg [7:0] \pageColumnIndex$next ;
  (* src = "sdram_controller.py:254" *)
  reg [14:0] powerUpCounter = 15'h0000;
  (* src = "sdram_controller.py:254" *)
  reg [14:0] \powerUpCounter$next ;
  (* enum_base_type = "SDRAMControllerStates" *)
  (* enum_value_000 = "InitOp" *)
  (* enum_value_001 = "ConfigurationOp" *)
  (* enum_value_010 = "Idle" *)
  (* enum_value_011 = "RefreshOp" *)
  (* enum_value_100 = "WriteBurstOp" *)
  (* enum_value_101 = "WriteOp" *)
  (* enum_value_110 = "ReadOp" *)
  (* enum_value_111 = "Error" *)
  (* src = "sdram_controller.py:227" *)
  reg [2:0] previousControllerState = 3'h0;
  (* src = "sdram_controller.py:227" *)
  reg [2:0] \previousControllerState$next ;
  (* src = "sdram_controller.py:252" *)
  reg refreshCmdIndex = 1'h0;
  (* src = "sdram_controller.py:252" *)
  reg \refreshCmdIndex$next ;
  (* src = "sdram_controller.py:253" *)
  reg refreshRequired = 1'h0;
  (* src = "sdram_controller.py:253" *)
  reg \refreshRequired$next ;
  (* src = "sdram_controller.py:702" *)
  reg repeatRefresh = 1'h0;
  (* src = "sdram_controller.py:702" *)
  reg \repeatRefresh$next ;
  (* src = "sdram_controller.py:201" *)
  output [10:0] sdramAddress;
  reg [10:0] sdramAddress = 11'h000;
  (* src = "sdram_controller.py:201" *)
  reg [10:0] \sdramAddress$next ;
  (* src = "sdram_controller.py:202" *)
  output [1:0] sdramBank;
  reg [1:0] sdramBank = 2'h0;
  (* src = "sdram_controller.py:202" *)
  reg [1:0] \sdramBank$next ;
  (* src = "sdram_controller.py:198" *)
  output sdramCASn;
  reg sdramCASn = 1'h0;
  (* src = "sdram_controller.py:198" *)
  reg \sdramCASn$next ;
  (* src = "sdram_controller.py:200" *)
  output sdramCSn;
  reg sdramCSn = 1'h0;
  (* src = "sdram_controller.py:200" *)
  reg \sdramCSn$next ;
  (* src = "sdram_controller.py:195" *)
  output sdramClk;
  wire sdramClk;
  (* src = "sdram_controller.py:196" *)
  output sdramClkEn;
  reg sdramClkEn = 1'h0;
  (* src = "sdram_controller.py:196" *)
  reg \sdramClkEn$next ;
  (* src = "sdram_controller.py:704" *)
  reg [2:0] sdramCtrlr_state = 3'h0;
  (* src = "sdram_controller.py:704" *)
  reg [2:0] \sdramCtrlr_state$next ;
  (* src = "sdram_controller.py:206" *)
  output [3:0] sdramDataMasks;
  reg [3:0] sdramDataMasks = 4'hf;
  (* src = "sdram_controller.py:206" *)
  reg [3:0] \sdramDataMasks$next ;
  (* src = "sdram_controller.py:204" *)
  output [31:0] sdramDqIn;
  reg [31:0] sdramDqIn = 32'd0;
  (* src = "sdram_controller.py:204" *)
  reg [31:0] \sdramDqIn$next ;
  (* src = "sdram_controller.py:203" *)
  input [31:0] sdramDqOut;
  wire [31:0] sdramDqOut;
  (* src = "sdram_controller.py:205" *)
  output sdramDqWRn;
  reg sdramDqWRn = 1'h0;
  (* src = "sdram_controller.py:205" *)
  reg \sdramDqWRn$next ;
  (* src = "sdram_controller.py:197" *)
  output sdramRASn;
  reg sdramRASn = 1'h0;
  (* src = "sdram_controller.py:197" *)
  reg \sdramRASn$next ;
  (* src = "sdram_controller.py:199" *)
  output sdramWEn;
  reg sdramWEn = 1'h0;
  (* src = "sdram_controller.py:199" *)
  reg \sdramWEn$next ;
  (* src = "sdram_controller.py:229" *)
  wire [1:0] targetBankAddress;
  (* src = "sdram_controller.py:236" *)
  reg targetBankCanActivate = 1'h0;
  (* src = "sdram_controller.py:236" *)
  reg \targetBankCanActivate$next ;
  (* src = "sdram_controller.py:237" *)
  reg targetBankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:237" *)
  reg \targetBankCanPreCharge$next ;
  (* src = "sdram_controller.py:238" *)
  reg [9:0] targetBankRefreshCounter = 10'h000;
  (* src = "sdram_controller.py:238" *)
  reg [9:0] \targetBankRefreshCounter$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:239" *)
  reg [2:0] targetBankState;
  (* src = "sdram_controller.py:231" *)
  wire [7:0] targetColumnAddress;
  (* src = "sdram_controller.py:232" *)
  wire [3:0] targetMask;
  (* src = "sdram_controller.py:230" *)
  wire [10:0] targetRowAddress;
  assign \$9  = cmdIndex == (* src = "sdram_controller.py:722" *) 1'h1;
  assign \$99  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$1000  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$1002  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1006  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1008  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$1012  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1014  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$101  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1020  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1022  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1024  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1026  = \$1022  | (* src = "sdram_controller.py:325" *) \$1024 ;
  assign \$1028  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1032  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1034  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1036  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$1038  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$103  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1040  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$1042  = \$1038  & (* src = "sdram_controller.py:439" *) \$1040 ;
  assign \$1046  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$1050  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1052  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1054  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1056  = \$1052  | (* src = "sdram_controller.py:325" *) \$1054 ;
  assign \$1058  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$105  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$1062  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$1066  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1068  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1070  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$1072  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$1074  = \$1070  & (* src = "sdram_controller.py:395" *) \$1072 ;
  assign \$1078  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$107  = ! (* src = "sdram_controller.py:1020" *) pageColumnIndex;
  assign \$1080  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1084  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1086  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1090  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$1092  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1096  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1098  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$109  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$1102  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1104  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1110  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1112  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1114  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1116  = \$1112  | (* src = "sdram_controller.py:325" *) \$1114 ;
  assign \$1118  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$111  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$1122  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1124  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1126  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$1128  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$1130  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$1132  = \$1128  & (* src = "sdram_controller.py:439" *) \$1130 ;
  assign \$1136  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$113  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1140  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1142  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1144  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1146  = \$1142  | (* src = "sdram_controller.py:325" *) \$1144 ;
  assign \$1148  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1152  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$1156  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1158  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$115  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1160  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$1162  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$1164  = \$1160  & (* src = "sdram_controller.py:395" *) \$1162 ;
  assign \$1168  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1170  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1174  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1176  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$117  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$1180  = cmdIndex == (* src = "sdram_controller.py:722" *) 1'h1;
  assign \$1182  = powerUpCounter > (* src = "sdram_controller.py:723" *) 1'h0;
  assign \$1184  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1188  = $signed(delayCounter) > (* src = "sdram_controller.py:386" *) $signed(4'h0);
  assign \$1190  = ! (* src = "sdram_controller.py:388" *) $signed(delayCounter);
  assign \$1193  = $signed(delayCounter) - (* src = "sdram_controller.py:387" *) $signed(4'h1);
  assign \$1195  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1197  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$11  = powerUpCounter > (* src = "sdram_controller.py:723" *) 1'h0;
  assign \$119  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1201  = $signed(delayCounter) > (* src = "sdram_controller.py:497" *) $signed(4'h0);
  assign \$1203  = ! (* src = "sdram_controller.py:499" *) $signed(delayCounter);
  assign \$1206  = $signed(delayCounter) - (* src = "sdram_controller.py:498" *) $signed(4'h1);
  assign \$1208  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$1210  = cmdIndex == (* src = "sdram_controller.py:763" *) 3'h5;
  assign \$1212  = $signed(delayCounter) > (* src = "sdram_controller.py:764" *) $signed(4'h0);
  assign \$1214  = ! (* src = "sdram_controller.py:766" *) $signed(delayCounter);
  assign \$1217  = $signed(delayCounter) - (* src = "sdram_controller.py:765" *) $signed(4'h1);
  assign \$1219  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$1221  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1223  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1225  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$1228  = $signed(delayCounter) - (* src = "sdram_controller.py:839" *) $signed(4'h1);
  assign \$1230  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$1232  = cmdIndex == (* src = "sdram_controller.py:932" *) 4'ha;
  assign \$1234  = $signed(delayCounter) > (* src = "sdram_controller.py:934" *) $signed(4'h0);
  assign \$1237  = $signed(delayCounter) - (* src = "sdram_controller.py:935" *) $signed(4'h1);
  assign \$123  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$1239  = ! (* src = "sdram_controller.py:936" *) $signed(delayCounter);
  assign \$1241  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$1243  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1245  = $signed(delayCounter) > (* src = "sdram_controller.py:997" *) $signed(4'h0);
  assign \$1248  = $signed(delayCounter) - (* src = "sdram_controller.py:998" *) $signed(4'h1);
  assign \$1250  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1252  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$1254  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$1256  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$1258  = $signed(delayCounter) > (* src = "sdram_controller.py:1065" *) $signed(4'h0);
  assign \$125  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1261  = $signed(delayCounter) - (* src = "sdram_controller.py:1066" *) $signed(4'h1);
  assign \$1263  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1265  = $signed(delayCounter) > (* src = "sdram_controller.py:1070" *) $signed(4'h0);
  assign \$1268  = $signed(delayCounter) - (* src = "sdram_controller.py:1071" *) $signed(4'h1);
  assign \$1270  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1272  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$1274  = $signed(delayCounter) > (* src = "sdram_controller.py:1080" *) $signed(4'h0);
  assign \$1277  = $signed(delayCounter) - (* src = "sdram_controller.py:1081" *) $signed(4'h1);
  assign \$127  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$1279  = ! (* src = "sdram_controller.py:1082" *) $signed(delayCounter);
  assign \$1281  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1285  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$1287  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$1289  = \$1287  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$1292  = $signed(delayCounter) - (* src = "sdram_controller.py:1102" *) $signed(4'h1);
  assign \$1294  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1298  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$129  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1300  = ! (* src = "sdram_controller.py:748" *) cmdRemainingCyclesCounter;
  assign \$1302  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1304  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1306  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1308  = \$1304  | (* src = "sdram_controller.py:325" *) \$1306 ;
  assign \$1310  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1314  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1316  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1318  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$131  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1320  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$1322  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$1324  = \$1320  & (* src = "sdram_controller.py:439" *) \$1322 ;
  assign \$1328  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$1332  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1334  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1336  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1338  = \$1334  | (* src = "sdram_controller.py:325" *) \$1336 ;
  assign \$133  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$1340  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1344  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1346  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1348  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$1350  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$1352  = \$1348  & (* src = "sdram_controller.py:395" *) \$1350 ;
  assign \$1356  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1358  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$135  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1362  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1366  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1368  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1372  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$1374  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1376  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1378  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$137  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$1380  = \$1376  | (* src = "sdram_controller.py:325" *) \$1378 ;
  assign \$1382  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1386  = ! (* src = "sdram_controller.py:334" *) targetBankAddress;
  assign \$1388  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$1392  = ! (* src = "sdram_controller.py:359" *) targetBankAddress;
  assign \$1394  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1396  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1398  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$13  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$139  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1400  = \$1396  | (* src = "sdram_controller.py:325" *) \$1398 ;
  assign \$1402  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1406  = ! (* src = "sdram_controller.py:334" *) targetBankAddress;
  assign \$1408  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1410  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1414  = ! (* src = "sdram_controller.py:359" *) targetBankAddress;
  assign \$1416  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1418  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$141  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1424  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$1426  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$1428  = \$1426  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$1430  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1434  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1436  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$143  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$1440  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$1442  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1444  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1446  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1448  = \$1444  | (* src = "sdram_controller.py:325" *) \$1446 ;
  assign \$1450  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1454  = targetBankAddress == (* src = "sdram_controller.py:334" *) 1'h1;
  assign \$1456  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$145  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$1460  = targetBankAddress == (* src = "sdram_controller.py:359" *) 1'h1;
  assign \$1462  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1464  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1466  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1468  = \$1464  | (* src = "sdram_controller.py:325" *) \$1466 ;
  assign \$1470  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1474  = targetBankAddress == (* src = "sdram_controller.py:334" *) 1'h1;
  assign \$1476  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1478  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$147  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$1482  = targetBankAddress == (* src = "sdram_controller.py:359" *) 1'h1;
  assign \$1484  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1486  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1492  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$1494  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$1496  = \$1494  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$1498  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$149  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$1502  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1504  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1508  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$1510  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1512  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1514  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1516  = \$1512  | (* src = "sdram_controller.py:325" *) \$1514 ;
  assign \$1518  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$151  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$1522  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h2;
  assign \$1524  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$1528  = targetBankAddress == (* src = "sdram_controller.py:359" *) 2'h2;
  assign \$1530  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1532  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1534  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1536  = \$1532  | (* src = "sdram_controller.py:325" *) \$1534 ;
  assign \$1538  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$153  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$1542  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h2;
  assign \$1544  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1546  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1550  = targetBankAddress == (* src = "sdram_controller.py:359" *) 2'h2;
  assign \$1552  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1554  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$155  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1560  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$1562  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$1564  = \$1562  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$1566  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1570  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$1572  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1576  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$1578  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$157  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$1580  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1582  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1584  = \$1580  | (* src = "sdram_controller.py:325" *) \$1582 ;
  assign \$1586  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1590  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h3;
  assign \$1592  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$1596  = targetBankAddress == (* src = "sdram_controller.py:359" *) 2'h3;
  assign \$1598  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$15  = ctrlWr & (* src = "sdram_controller.py:797" *) burstWritesMode;
  assign \$159  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1600  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1602  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1604  = \$1600  | (* src = "sdram_controller.py:325" *) \$1602 ;
  assign \$1606  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1610  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h3;
  assign \$1612  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1614  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1618  = targetBankAddress == (* src = "sdram_controller.py:359" *) 2'h3;
  assign \$161  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1620  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1622  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1628  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$1630  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$1632  = \$1630  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$1634  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1636  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$1638  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$163  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$1640  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1642  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1644  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1646  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1648  = \$1644  | (* src = "sdram_controller.py:325" *) \$1646 ;
  assign \$1650  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1654  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1656  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1658  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$165  = ! (* src = "sdram_controller.py:1020" *) pageColumnIndex;
  assign \$1660  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$1662  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$1664  = \$1660  & (* src = "sdram_controller.py:439" *) \$1662 ;
  assign \$1666  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$1668  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$1670  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$1672  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$1674  = \$1670  & (* src = "sdram_controller.py:609" *) \$1672 ;
  assign \$1676  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1678  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$167  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$1680  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1682  = \$1678  | (* src = "sdram_controller.py:325" *) \$1680 ;
  assign \$1684  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1688  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1690  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1692  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$1694  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$1696  = \$1692  & (* src = "sdram_controller.py:395" *) \$1694 ;
  assign \$1698  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$169  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$1700  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$1702  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$1704  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$1706  = \$1702  & (* src = "sdram_controller.py:609" *) \$1704 ;
  assign \$1708  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1710  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$1712  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1714  = ! (* src = "sdram_controller.py:748" *) cmdRemainingCyclesCounter;
  assign \$1716  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1718  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$171  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$1720  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1722  = \$1718  | (* src = "sdram_controller.py:325" *) \$1720 ;
  assign \$1724  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1728  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$1730  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$1732  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$1734  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$1736  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$1738  = \$1734  & (* src = "sdram_controller.py:439" *) \$1736 ;
  assign \$173  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$1742  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1744  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1746  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1748  = \$1744  | (* src = "sdram_controller.py:325" *) \$1746 ;
  assign \$1750  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1754  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$1756  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$1758  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$175  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$1760  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$1762  = \$1758  & (* src = "sdram_controller.py:395" *) \$1760 ;
  assign \$1766  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1768  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$1770  = ctrlWr & (* src = "sdram_controller.py:797" *) burstWritesMode;
  assign \$1772  = cmdIndex == (* src = "sdram_controller.py:932" *) 4'ha;
  assign \$1774  = ! (* src = "sdram_controller.py:936" *) $signed(delayCounter);
  assign \$1776  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$1778  = ! (* src = "sdram_controller.py:1082" *) $signed(delayCounter);
  assign \$177  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$1780  = ctrlWr & (* src = "sdram_controller.py:797" *) burstWritesMode;
  assign \$1782  = ! (* src = "sdram_controller.py:814" *) cmdIndex;
  assign \$1784  = 9'h100 - (* src = "sdram_controller.py:818" *) targetColumnAddress;
  assign \$1788  = \$1786  + (* src = "sdram_controller.py:818" *) 4'hf;
  assign \$1790  = \$1788  + (* src = "sdram_controller.py:818" *) 3'h5;
  assign \$1792  = targetBankRefreshCounter < (* src = "sdram_controller.py:818" *) \$1790 ;
  assign \$1794  = ! (* src = "sdram_controller.py:951" *) cmdIndex;
  assign \$1796  = 9'h100 - (* src = "sdram_controller.py:953" *) targetColumnAddress;
  assign \$17  = ~ (* src = "sdram_controller.py:795" *) ctrlReady;
  assign \$1800  = \$1798  + (* src = "sdram_controller.py:953" *) 4'hd;
  assign \$1802  = \$1800  + (* src = "sdram_controller.py:953" *) 3'h5;
  assign \$1804  = targetBankRefreshCounter < (* src = "sdram_controller.py:953" *) \$1802 ;
  assign \$1808  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$1810  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$1812  = \$1810  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$1814  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1816  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1818  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$181  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$1820  = \$1816  | (* src = "sdram_controller.py:325" *) \$1818 ;
  assign \$1822  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1826  = ! (* src = "sdram_controller.py:334" *) targetBankAddress;
  assign \$1828  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1830  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1832  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1834  = \$1830  | (* src = "sdram_controller.py:325" *) \$1832 ;
  assign \$1836  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$183  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$1840  = ! (* src = "sdram_controller.py:334" *) targetBankAddress;
  assign \$1842  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1844  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1846  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1848  = \$1844  | (* src = "sdram_controller.py:325" *) \$1846 ;
  assign \$1850  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1854  = ! (* src = "sdram_controller.py:334" *) targetBankAddress;
  assign \$1856  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1858  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$185  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$1860  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1862  = \$1858  | (* src = "sdram_controller.py:325" *) \$1860 ;
  assign \$1864  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1868  = ! (* src = "sdram_controller.py:334" *) targetBankAddress;
  assign \$1870  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1872  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1874  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1876  = \$1872  | (* src = "sdram_controller.py:325" *) \$1874 ;
  assign \$1878  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$187  = ~ (* src = "sdram_controller.py:371" *) sdramClkEn;
  assign \$1882  = targetBankAddress == (* src = "sdram_controller.py:334" *) 1'h1;
  assign \$1884  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1886  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1888  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1890  = \$1886  | (* src = "sdram_controller.py:325" *) \$1888 ;
  assign \$1892  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1896  = targetBankAddress == (* src = "sdram_controller.py:334" *) 1'h1;
  assign \$1898  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$189  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$1900  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1902  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1904  = \$1900  | (* src = "sdram_controller.py:325" *) \$1902 ;
  assign \$1906  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1910  = targetBankAddress == (* src = "sdram_controller.py:334" *) 1'h1;
  assign \$1912  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1914  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1916  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1918  = \$1914  | (* src = "sdram_controller.py:325" *) \$1916 ;
  assign \$191  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$1920  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1924  = targetBankAddress == (* src = "sdram_controller.py:334" *) 1'h1;
  assign \$1926  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1928  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1930  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1932  = \$1928  | (* src = "sdram_controller.py:325" *) \$1930 ;
  assign \$1934  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1938  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h2;
  assign \$193  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$1940  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1942  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1944  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1946  = \$1942  | (* src = "sdram_controller.py:325" *) \$1944 ;
  assign \$1948  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1952  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h2;
  assign \$1954  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1956  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1958  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$195  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$1960  = \$1956  | (* src = "sdram_controller.py:325" *) \$1958 ;
  assign \$1962  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1966  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h2;
  assign \$1968  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1970  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1972  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1974  = \$1970  | (* src = "sdram_controller.py:325" *) \$1972 ;
  assign \$1976  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$197  = ~ (* src = "sdram_controller.py:486" *) sdramClkEn;
  assign \$1980  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h2;
  assign \$1982  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$1984  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1986  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$1988  = \$1984  | (* src = "sdram_controller.py:325" *) \$1986 ;
  assign \$1990  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$1994  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h3;
  assign \$1996  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$1998  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$1  = bankController0_bankState != (* src = "sdram_controller.py:655" *) 1'h1;
  assign \$19  = ~ (* src = "sdram_controller.py:801" *) ctrlReady;
  assign \$199  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$2000  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$2002  = \$1998  | (* src = "sdram_controller.py:325" *) \$2000 ;
  assign \$2004  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$2008  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h3;
  assign \$2010  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$2012  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$2014  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$2016  = \$2012  | (* src = "sdram_controller.py:325" *) \$2014 ;
  assign \$2018  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$201  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$2022  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h3;
  assign \$2024  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$2026  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$2028  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$2030  = \$2026  | (* src = "sdram_controller.py:325" *) \$2028 ;
  assign \$2032  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$2036  = targetBankAddress == (* src = "sdram_controller.py:334" *) 2'h3;
  assign \$2038  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$203  = ~ (* src = "sdram_controller.py:546" *) sdramClkEn;
  assign \$2040  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$2042  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$2044  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$2046  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$2048  = \$2044  & (* src = "sdram_controller.py:609" *) \$2046 ;
  assign \$2052  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$2054  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$2056  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$2058  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$2060  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$2062  = \$2058  & (* src = "sdram_controller.py:395" *) \$2060 ;
  assign \$2066  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$2068  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$2070  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$2072  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$2074  = \$2070  & (* src = "sdram_controller.py:609" *) \$2072 ;
  assign \$2078  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$207  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$2080  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$2082  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$2084  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$2086  = pageColumnIndex < (* src = "sdram_controller.py:910" *) 8'hff;
  assign \$2089  = pageColumnIndex + (* src = "sdram_controller.py:911" *) 1'h1;
  assign \$2091  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$2093  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$2095  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$2097  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$209  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$2100  = pageColumnIndex + (* src = "sdram_controller.py:1053" *) 1'h1;
  assign \$2102  = cmdIndex == (* src = "sdram_controller.py:862" *) 3'h6;
  assign \$2104  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$2106  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$2108  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$2110  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$2112  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$2114  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$2116  = $signed(delayCounter) > (* src = "sdram_controller.py:997" *) $signed(4'h0);
  assign \$2118  = $signed(delayCounter) == (* src = "sdram_controller.py:999" *) $signed(4'h2);
  assign \$211  = ~ (* src = "sdram_controller.py:505" *) sdramClkEn;
  assign \$2120  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$2122  = pageColumnIndex == (* src = "sdram_controller.py:1061" *) 8'hfc;
  assign \$2124  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$2126  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$2128  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$2130  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$2132  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$2134  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$2136  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$2138  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$213  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$2140  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$2142  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$2144  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$2146  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$2150  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$2152  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$2154  = \$2152  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  always @(posedge 1'h0)
    targetBankCanActivate <= \targetBankCanActivate$next ;
  always @(posedge 1'h0)
    targetBankCanPreCharge <= \targetBankCanPreCharge$next ;
  always @(posedge 1'h0)
    targetBankRefreshCounter <= \targetBankRefreshCounter$next ;
  always @(posedge 1'h0)
    sdramCtrlr_state <= \sdramCtrlr_state$next ;
  assign \$215  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  always @(posedge 1'h0)
    previousControllerState <= \previousControllerState$next ;
  always @(posedge 1'h0)
    currentCommand <= \currentCommand$next ;
  always @(posedge 1'h0)
    sdramClkEn <= \sdramClkEn$next ;
  always @(posedge 1'h0)
    sdramCSn <= \sdramCSn$next ;
  always @(posedge 1'h0)
    repeatRefresh <= \repeatRefresh$next ;
  always @(posedge 1'h0)
    powerUpCounter <= \powerUpCounter$next ;
  always @(posedge 1'h0)
    cmdIndex <= \cmdIndex$next ;
  always @(posedge 1'h0)
    sdramRASn <= \sdramRASn$next ;
  always @(posedge 1'h0)
    sdramCASn <= \sdramCASn$next ;
  always @(posedge 1'h0)
    sdramWEn <= \sdramWEn$next ;
  always @(posedge 1'h0)
    delayCounter <= \delayCounter$next ;
  always @(posedge 1'h0)
    sdramAddress <= \sdramAddress$next ;
  always @(posedge 1'h0)
    bankController0_bankState <= \bankController0_bankState$next ;
  always @(posedge 1'h0)
    bankController1_bankState <= \bankController1_bankState$next ;
  always @(posedge 1'h0)
    bankController2_bankState <= \bankController2_bankState$next ;
  always @(posedge 1'h0)
    bankController3_bankState <= \bankController3_bankState$next ;
  always @(posedge 1'h0)
    errorState <= \errorState$next ;
  always @(posedge 1'h0)
    sdramBank <= \sdramBank$next ;
  always @(posedge 1'h0)
    burstWritesMode <= \burstWritesMode$next ;
  always @(posedge 1'h0)
    ctrlReady <= \ctrlReady$next ;
  assign \$217  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  always @(posedge 1'h0)
    ctrlAddress <= \ctrlAddress$next ;
  always @(posedge 1'h0)
    refreshRequired <= \refreshRequired$next ;
  always @(posedge 1'h0)
    sdramDataMasks <= \sdramDataMasks$next ;
  always @(posedge 1'h0)
    pageColumnIndex <= \pageColumnIndex$next ;
  always @(posedge 1'h0)
    ctrlRdInProgress <= \ctrlRdInProgress$next ;
  always @(posedge 1'h0)
    ctrlRdIncAddress <= \ctrlRdIncAddress$next ;
  always @(posedge 1'h0)
    ctrlWrIncAddress <= \ctrlWrIncAddress$next ;
  always @(posedge 1'h0)
    sdramDqWRn <= \sdramDqWRn$next ;
  always @(posedge 1'h0)
    sdramDqIn <= \sdramDqIn$next ;
  always @(posedge 1'h0)
    ctrlWrInProgress <= \ctrlWrInProgress$next ;
  always @(posedge 1'h0)
    refreshCmdIndex <= \refreshCmdIndex$next ;
  assign \$21  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$219  = \$215  | (* src = "sdram_controller.py:325" *) \$217 ;
  assign \$221  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$225  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$227  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$229  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$231  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$233  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$235  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$237  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$23  = cmdIndex == (* src = "sdram_controller.py:932" *) 4'ha;
  assign \$239  = \$235  & (* src = "sdram_controller.py:439" *) \$237 ;
  assign \$241  = ~ (* src = "sdram_controller.py:443" *) sdramClkEn;
  assign \$243  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$245  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$247  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$249  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$251  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$253  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$255  = \$251  & (* src = "sdram_controller.py:609" *) \$253 ;
  assign \$257  = ~ (* src = "sdram_controller.py:613" *) sdramClkEn;
  assign \$25  = ! (* src = "sdram_controller.py:936" *) $signed(delayCounter);
  assign \$259  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$261  = ~ (* src = "sdram_controller.py:352" *) sdramClkEn;
  assign \$263  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$265  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$267  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$269  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$271  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$273  = \$269  | (* src = "sdram_controller.py:325" *) \$271 ;
  assign \$275  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$27  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$279  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$281  = ~ (* src = "sdram_controller.py:505" *) sdramClkEn;
  assign \$283  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$285  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$287  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$289  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$291  = \$287  & (* src = "sdram_controller.py:395" *) \$289 ;
  assign \$293  = ~ (* src = "sdram_controller.py:399" *) sdramClkEn;
  assign \$295  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$297  = ! (* src = "sdram_controller.py:1020" *) pageColumnIndex;
  assign \$29  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$299  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$301  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$303  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$305  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$307  = \$303  & (* src = "sdram_controller.py:609" *) \$305 ;
  assign \$309  = ~ (* src = "sdram_controller.py:613" *) sdramClkEn;
  assign \$311  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$313  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$315  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$317  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$31  = ! (* src = "sdram_controller.py:1082" *) $signed(delayCounter);
  assign \$319  = ~ (* src = "sdram_controller.py:352" *) sdramClkEn;
  assign \$321  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$323  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$325  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$327  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$329  = ~ (* src = "sdram_controller.py:546" *) sdramClkEn;
  assign \$335  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$337  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$339  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$343  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$345  = ~ (* src = "sdram_controller.py:371" *) sdramClkEn;
  assign \$349  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$351  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$355  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$357  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$35  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$359  = ~ (* src = "sdram_controller.py:486" *) sdramClkEn;
  assign \$363  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$365  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$367  = ~ (* src = "sdram_controller.py:546" *) sdramClkEn;
  assign \$371  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$373  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$377  = ~ (* src = "sdram_controller.py:505" *) sdramClkEn;
  assign \$37  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$381  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$383  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$385  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$387  = \$383  | (* src = "sdram_controller.py:325" *) \$385 ;
  assign \$389  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$393  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$395  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$3  = bankController1_bankState != (* src = "sdram_controller.py:655" *) 1'h1;
  assign \$39  = \$37  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$399  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$401  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$403  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$405  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$407  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$409  = \$405  & (* src = "sdram_controller.py:439" *) \$407 ;
  assign \$411  = ~ (* src = "sdram_controller.py:443" *) sdramClkEn;
  assign \$415  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$417  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$41  = previousControllerState == (* src = "sdram_controller.py:1110" *) 3'h4;
  assign \$421  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$423  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$425  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$427  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$429  = \$425  & (* src = "sdram_controller.py:609" *) \$427 ;
  assign \$431  = ~ (* src = "sdram_controller.py:613" *) sdramClkEn;
  assign \$435  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$437  = ~ (* src = "sdram_controller.py:352" *) sdramClkEn;
  assign \$43  = previousControllerState == (* src = "sdram_controller.py:1112" *) 3'h6;
  assign \$441  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$443  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$447  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$449  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$451  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$453  = \$449  | (* src = "sdram_controller.py:325" *) \$451 ;
  assign \$455  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$45  = cmdIndex == (* src = "sdram_controller.py:722" *) 1'h1;
  assign \$459  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$461  = ~ (* src = "sdram_controller.py:505" *) sdramClkEn;
  assign \$465  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$467  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$469  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$471  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$473  = \$469  & (* src = "sdram_controller.py:395" *) \$471 ;
  assign \$475  = ~ (* src = "sdram_controller.py:399" *) sdramClkEn;
  assign \$47  = powerUpCounter > (* src = "sdram_controller.py:723" *) 1'h0;
  assign \$479  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$481  = ! (* src = "sdram_controller.py:1020" *) pageColumnIndex;
  assign \$483  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$487  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$489  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$491  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$493  = \$489  & (* src = "sdram_controller.py:609" *) \$491 ;
  assign \$495  = ~ (* src = "sdram_controller.py:613" *) sdramClkEn;
  assign \$49  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$499  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$501  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$505  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$507  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$509  = ~ (* src = "sdram_controller.py:352" *) sdramClkEn;
  assign \$513  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$515  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$51  = ctrlWr & (* src = "sdram_controller.py:797" *) burstWritesMode;
  assign \$519  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$521  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$523  = ~ (* src = "sdram_controller.py:546" *) sdramClkEn;
  assign \$529  = ~ (* src = "sdram_controller.py:533" *) sdramClkEn;
  assign \$533  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$537  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$53  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$539  = $signed(delayCounter) > (* src = "sdram_controller.py:386" *) $signed(4'h0);
  assign \$541  = ! (* src = "sdram_controller.py:388" *) $signed(delayCounter);
  assign \$543  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$547  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$549  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$551  = $signed(delayCounter) > (* src = "sdram_controller.py:497" *) $signed(4'h0);
  assign \$553  = ! (* src = "sdram_controller.py:499" *) $signed(delayCounter);
  assign \$555  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$557  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$55  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$561  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$567  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$569  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$571  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$573  = \$569  | (* src = "sdram_controller.py:325" *) \$571 ;
  assign \$575  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$579  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$583  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$585  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$587  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$589  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$591  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$593  = \$589  & (* src = "sdram_controller.py:439" *) \$591 ;
  assign \$597  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$5  = bankController2_bankState != (* src = "sdram_controller.py:655" *) 1'h1;
  assign \$59  = $signed(delayCounter) > (* src = "sdram_controller.py:1101" *) $signed(4'h0);
  assign \$601  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$603  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$605  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$607  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$609  = \$605  & (* src = "sdram_controller.py:609" *) \$607 ;
  assign \$613  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$617  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$61  = ! (* src = "sdram_controller.py:1103" *) $signed(delayCounter);
  assign \$621  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$623  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$625  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$627  = \$623  | (* src = "sdram_controller.py:325" *) \$625 ;
  assign \$629  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$633  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$637  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$63  = \$61  & (* src = "sdram_controller.py:1103" *) cmdCompleted;
  assign \$639  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$641  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$643  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$645  = \$641  & (* src = "sdram_controller.py:395" *) \$643 ;
  assign \$649  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$651  = ! (* src = "sdram_controller.py:1020" *) pageColumnIndex;
  assign \$655  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$657  = targetBankState != (* src = "sdram_controller.py:609" *) 2'h2;
  assign \$65  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$659  = targetBankState != (* src = "sdram_controller.py:610" *) 2'h3;
  assign \$661  = \$657  & (* src = "sdram_controller.py:609" *) \$659 ;
  assign \$665  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$669  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$671  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$675  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$67  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$679  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$681  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$689  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$693  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$697  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$69  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$701  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$703  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$707  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$709  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$713  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$71  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$719  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$721  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$723  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$725  = \$721  | (* src = "sdram_controller.py:325" *) \$723 ;
  assign \$727  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$731  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$735  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$737  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$73  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$739  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$741  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$743  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$745  = \$741  & (* src = "sdram_controller.py:439" *) \$743 ;
  assign \$749  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$753  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$757  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$75  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$761  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$763  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$765  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$767  = \$763  | (* src = "sdram_controller.py:325" *) \$765 ;
  assign \$769  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$773  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$777  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$77  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$779  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$781  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$783  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$785  = \$781  & (* src = "sdram_controller.py:395" *) \$783 ;
  assign \$789  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$791  = ! (* src = "sdram_controller.py:1020" *) pageColumnIndex;
  assign \$795  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$7  = bankController3_bankState != (* src = "sdram_controller.py:655" *) 1'h1;
  assign \$79  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$799  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$801  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$805  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$809  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$811  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$81  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$819  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$821  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$823  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$825  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$827  = cmdIndex == (* src = "sdram_controller.py:722" *) 1'h1;
  assign \$829  = powerUpCounter > (* src = "sdram_controller.py:723" *) 1'h0;
  assign \$832  = powerUpCounter - (* src = "sdram_controller.py:724" *) 1'h1;
  assign \$834  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$836  = cmdIndex == (* src = "sdram_controller.py:722" *) 1'h1;
  assign \$838  = powerUpCounter > (* src = "sdram_controller.py:723" *) 1'h0;
  assign \$83  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$840  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$842  = cmdIndex == (* src = "sdram_controller.py:742" *) 1'h1;
  assign \$844  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$846  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$848  = cmdIndex == (* src = "sdram_controller.py:758" *) 3'h4;
  assign \$850  = cmdIndex == (* src = "sdram_controller.py:763" *) 3'h5;
  assign \$852  = $signed(delayCounter) > (* src = "sdram_controller.py:764" *) $signed(4'h0);
  assign \$854  = ! (* src = "sdram_controller.py:766" *) $signed(delayCounter);
  assign \$856  = cmdIndex == (* src = "sdram_controller.py:769" *) 3'h6;
  assign \$858  = ! (* src = "sdram_controller.py:814" *) cmdIndex;
  assign \$85  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$860  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$862  = cmdIndex == (* src = "sdram_controller.py:831" *) 2'h2;
  assign \$864  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$866  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$868  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$870  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$872  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h5;
  assign \$874  = cmdIndex == (* src = "sdram_controller.py:862" *) 3'h6;
  assign \$876  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$878  = pageColumnIndex < (* src = "sdram_controller.py:910" *) 8'hff;
  assign \$87  = cmdIndex == (* src = "sdram_controller.py:849" *) 3'h4;
  assign \$880  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$882  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$884  = cmdIndex == (* src = "sdram_controller.py:932" *) 4'ha;
  assign \$886  = ! (* src = "sdram_controller.py:936" *) $signed(delayCounter);
  assign \$888  = ! (* src = "sdram_controller.py:951" *) cmdIndex;
  assign \$890  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$892  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$894  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$896  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$898  = cmdIndex == (* src = "sdram_controller.py:1013" *) 3'h4;
  assign \$89  = cmdIndex == (* src = "sdram_controller.py:869" *) 3'h7;
  assign \$900  = pageColumnIndex < (* src = "sdram_controller.py:1052" *) 8'hff;
  assign \$902  = cmdIndex == (* src = "sdram_controller.py:1063" *) 3'h5;
  assign \$904  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$906  = cmdIndex == (* src = "sdram_controller.py:1078" *) 3'h7;
  assign \$908  = ! (* src = "sdram_controller.py:1082" *) $signed(delayCounter);
  assign \$910  = ! (* src = "sdram_controller.py:712" *) cmdIndex;
  assign \$912  = ! (* src = "sdram_controller.py:737" *) cmdIndex;
  assign \$916  = cmdIndex == (* src = "sdram_controller.py:746" *) 2'h2;
  assign \$918  = ~ (* src = "sdram_controller.py:483" *) allBanksIdle;
  assign \$91  = pageColumnIndex == (* src = "sdram_controller.py:915" *) 8'hfe;
  assign \$922  = cmdIndex == (* src = "sdram_controller.py:754" *) 2'h3;
  assign \$924  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  assign \$930  = cmdIndex == (* src = "sdram_controller.py:820" *) 1'h1;
  assign \$932  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$934  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$936  = \$932  | (* src = "sdram_controller.py:325" *) \$934 ;
  assign \$938  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$93  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$942  = cmdIndex == (* src = "sdram_controller.py:837" *) 2'h3;
  assign \$944  = $signed(delayCounter) > (* src = "sdram_controller.py:838" *) $signed(4'h0);
  assign \$946  = ! (* src = "sdram_controller.py:840" *) $signed(delayCounter);
  assign \$948  = targetBankState != (* src = "sdram_controller.py:439" *) 2'h2;
  assign \$950  = targetBankState != (* src = "sdram_controller.py:440" *) 2'h3;
  assign \$952  = \$948  & (* src = "sdram_controller.py:439" *) \$950 ;
  assign \$956  = cmdIndex == (* src = "sdram_controller.py:917" *) 4'h8;
  assign \$95  = cmdIndex == (* src = "sdram_controller.py:926" *) 4'h9;
  assign \$960  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$962  = targetBankState != (* src = "sdram_controller.py:325" *) 1'h1;
  assign \$964  = ~ (* src = "sdram_controller.py:325" *) targetBankCanActivate;
  assign \$966  = \$962  | (* src = "sdram_controller.py:325" *) \$964 ;
  assign \$968  = ~ (* src = "sdram_controller.py:327" *) sdramClkEn;
  assign \$972  = cmdIndex == (* src = "sdram_controller.py:965" *) 2'h2;
  assign \$976  = cmdIndex == (* src = "sdram_controller.py:970" *) 2'h3;
  assign \$978  = ! (* src = "sdram_controller.py:1001" *) $signed(delayCounter);
  assign \$97  = cmdIndex == (* src = "sdram_controller.py:955" *) 1'h1;
  assign \$980  = targetBankState != (* src = "sdram_controller.py:395" *) 2'h2;
  assign \$982  = targetBankState != (* src = "sdram_controller.py:396" *) 2'h3;
  assign \$984  = \$980  & (* src = "sdram_controller.py:395" *) \$982 ;
  assign \$988  = cmdIndex == (* src = "sdram_controller.py:1069" *) 3'h6;
  assign \$990  = ! (* src = "sdram_controller.py:1072" *) $signed(delayCounter);
  assign \$994  = ~ (* src = "sdram_controller.py:1094" *) refreshCmdIndex;
  assign \$996  = ~ (* src = "sdram_controller.py:543" *) allBanksIdle;
  bankController0 bankController0 (
    .bankActivated(bankController0_bankActivated),
    .bankCanActivate(bankController0_bankCanActivate),
    .bankCanPreCharge(bankController0_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController0_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController0_bankShouldRefresh),
    .bankState(bankController0_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController0_otherBankActivated)
  );
  bankController1 bankController1 (
    .bankActivated(bankController1_bankActivated),
    .bankCanActivate(bankController1_bankCanActivate),
    .bankCanPreCharge(bankController1_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController1_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController1_bankShouldRefresh),
    .bankState(bankController1_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController1_otherBankActivated)
  );
  bankController2 bankController2 (
    .bankActivated(bankController2_bankActivated),
    .bankCanActivate(bankController2_bankCanActivate),
    .bankCanPreCharge(bankController2_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController2_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController2_bankShouldRefresh),
    .bankState(bankController2_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController2_otherBankActivated)
  );
  bankController3 bankController3 (
    .bankActivated(bankController3_bankActivated),
    .bankCanActivate(bankController3_bankCanActivate),
    .bankCanPreCharge(bankController3_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController3_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController3_bankShouldRefresh),
    .bankState(bankController3_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController3_otherBankActivated)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    allBanksIdle = 1'h1;
    (* src = "sdram_controller.py:655" *)
    casez (\$1 )
      /* src = "sdram_controller.py:655" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
    (* src = "sdram_controller.py:655" *)
    casez (\$3 )
      /* src = "sdram_controller.py:655" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
    (* src = "sdram_controller.py:655" *)
    casez (\$5 )
      /* src = "sdram_controller.py:655" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
    (* src = "sdram_controller.py:655" *)
    casez (\$7 )
      /* src = "sdram_controller.py:655" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramCtrlr_state$next  = sdramCtrlr_state;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
        begin
          \sdramCtrlr_state$next  = 3'h0;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:722" *)
                casez (\$9 )
                  /* src = "sdram_controller.py:722" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:723" *)
                      casez (\$11 )
                        /* src = "sdram_controller.py:723" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:725" */
                        default:
                            \sdramCtrlr_state$next  = 3'h2;
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
        begin
          \sdramCtrlr_state$next  = 3'h2;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:736" */
            default:
                (* src = "sdram_controller.py:769" *)
                casez (\$13 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:772" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:772" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:775" */
                        default:
                            \sdramCtrlr_state$next  = 3'h3;
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
        begin
          \sdramCtrlr_state$next  = 3'h3;
          (* src = "sdram_controller.py:784" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:784" */
            2'b?1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:787" */
            2'b1?:
                (* src = "sdram_controller.py:788" *)
                casez ({ \$15 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:788" */
                  3'b??1:
                      \sdramCtrlr_state$next  = 3'h4;
                  /* src = "sdram_controller.py:791" */
                  3'b?1?:
                      (* src = "sdram_controller.py:795" *)
                      casez (\$17 )
                        /* src = "sdram_controller.py:795" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h5;
                      endcase
                  /* src = "sdram_controller.py:797" */
                  3'b1??:
                      (* src = "sdram_controller.py:801" *)
                      casez (\$19 )
                        /* src = "sdram_controller.py:801" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h6;
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
        begin
          \sdramCtrlr_state$next  = 3'h5;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$21 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            \sdramCtrlr_state$next  = 3'h4;
                      endcase
                endcase
                (* src = "sdram_controller.py:932" *)
                casez (\$23 )
                  /* src = "sdram_controller.py:932" */
                  1'h1:
                      (* src = "sdram_controller.py:936" *)
                      casez (\$25 )
                        /* src = "sdram_controller.py:936" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h3;
                      endcase
                endcase
              end
          endcase
        end
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
        begin
          \sdramCtrlr_state$next  = 3'h6;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$27 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            \sdramCtrlr_state$next  = 3'h4;
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$29 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      (* src = "sdram_controller.py:1082" *)
                      casez (\$31 )
                        /* src = "sdram_controller.py:1082" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h3;
                      endcase
                endcase
              end
          endcase
        end
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
        begin
          \sdramCtrlr_state$next  = 3'h4;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1099" *)
                casez (\$33 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$39 , \$35  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:1112" *)
                            casez (\$43 )
                              /* src = "sdram_controller.py:1112" */
                              1'h1:
                                  \sdramCtrlr_state$next  = 3'h5;
                              /* src = "sdram_controller.py:1114" */
                              default:
                                  \sdramCtrlr_state$next  = 3'h3;
                            endcase
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "Error/1" */
      /* src = "sdram_controller.py:1116" */
      3'h1:
          \sdramCtrlr_state$next  = 3'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramCtrlr_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    currentControllerState = 3'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          currentControllerState = 3'h0;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          currentControllerState = 3'h1;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          currentControllerState = 3'h2;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          currentControllerState = 3'h6;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          currentControllerState = 3'h4;
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          currentControllerState = 3'h3;
      /* \amaranth.decoding  = "Error/1" */
      /* src = "sdram_controller.py:1116" */
      3'h1:
          currentControllerState = 3'h7;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \previousControllerState$next  = previousControllerState;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:722" *)
                casez (\$45 )
                  /* src = "sdram_controller.py:722" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:723" *)
                      casez (\$47 )
                        /* src = "sdram_controller.py:723" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:725" */
                        default:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:736" */
            default:
                (* src = "sdram_controller.py:769" *)
                casez (\$49 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:772" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:772" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:775" */
                        default:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:784" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:784" */
            2'b?1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:787" */
            2'b1?:
                (* src = "sdram_controller.py:788" *)
                casez ({ \$51 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:788" */
                  3'b??1:
                      \previousControllerState$next  = currentControllerState;
                  /* src = "sdram_controller.py:791" */
                  3'b?1?:
                      \previousControllerState$next  = currentControllerState;
                  /* src = "sdram_controller.py:797" */
                  3'b1??:
                      \previousControllerState$next  = currentControllerState;
                endcase
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$53 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$55 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1099" *)
                casez (\$57 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$63 , \$59  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \previousControllerState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    nextCommand = 5'h00;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$65 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$67 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      nextCommand = 5'h03;
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$69 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$71 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      nextCommand = 5'h08;
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$73 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      nextCommand = 5'h0c;
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$75 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          nextCommand = 5'h09;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$77 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            nextCommand = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$79 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$81 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$85 , \$83  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            nextCommand = 5'h06;
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$87 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$89 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$91 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            nextCommand = 5'h12;
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$93 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            nextCommand = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$95 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$97 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            nextCommand = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$99 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      nextCommand = 5'h09;
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$101 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$103 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            nextCommand = 5'h04;
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$105 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1020" *)
                      casez (\$107 )
                        /* src = "sdram_controller.py:1020" */
                        1'h1:
                            nextCommand = 5'h0b;
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$109 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            nextCommand = 5'h12;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$111 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$113 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$115 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  nextCommand = 5'h02;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$117 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$119 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      nextCommand = 5'h0c;
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$121 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \currentCommand$next  = currentCommand;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$123 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$125 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      \currentCommand$next  = 5'h03;
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$127 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$129 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      \currentCommand$next  = 5'h08;
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$131 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      \currentCommand$next  = 5'h0c;
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$133 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          \currentCommand$next  = 5'h09;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$135 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            \currentCommand$next  = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$137 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$139 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$143 , \$141  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            \currentCommand$next  = 5'h06;
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$145 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$147 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$149 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            \currentCommand$next  = 5'h12;
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$151 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            \currentCommand$next  = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$153 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$155 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            \currentCommand$next  = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$157 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      \currentCommand$next  = 5'h09;
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$159 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$161 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            \currentCommand$next  = 5'h04;
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$163 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1020" *)
                      casez (\$165 )
                        /* src = "sdram_controller.py:1020" */
                        1'h1:
                            \currentCommand$next  = 5'h0b;
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$167 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            \currentCommand$next  = 5'h12;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$169 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$171 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$173 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  \currentCommand$next  = 5'h02;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$175 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$177 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      \currentCommand$next  = 5'h0c;
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$179 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \currentCommand$next  = 5'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramClkEn$next  = sdramClkEn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$181 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$183 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \sdramClkEn$next  = 1'h0;
                      endcase
                    end
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$185 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:371" *)
                      casez (\$187 )
                        /* src = "sdram_controller.py:371" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$189 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$191 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$193 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$195 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                            (* src = "sdram_controller.py:486" *)
                            casez (\$197 )
                              /* src = "sdram_controller.py:486" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$199 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$201 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                          begin
                            (* src = "sdram_controller.py:546" *)
                            casez (\$203 )
                              /* src = "sdram_controller.py:546" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                            (* src = "sdram_controller.py:549" *)
                            casez (\$205 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$207 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$209 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:505" *)
          casez (\$211 )
            /* src = "sdram_controller.py:505" */
            1'h1:
                \sdramClkEn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$213 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$223 , \$221 , \$219  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$225 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$227 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$229 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$233 , \$231  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$239 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:443" *)
                                  casez (\$241 )
                                    /* src = "sdram_controller.py:443" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$243 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$245 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$247 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$249 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$255 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                  (* src = "sdram_controller.py:613" *)
                                  casez (\$257 )
                                    /* src = "sdram_controller.py:613" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$259 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:352" *)
                            casez (\$261 )
                              /* src = "sdram_controller.py:352" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$263 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$265 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$267 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$277 , \$275 , \$273  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$279 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:505" *)
                      casez (\$281 )
                        /* src = "sdram_controller.py:505" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$283 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$285 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$291 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:399" *)
                                  casez (\$293 )
                                    /* src = "sdram_controller.py:399" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$295 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1020" *)
                      casez (\$297 )
                        /* src = "sdram_controller.py:1020" */
                        1'h1:
                            (* src = "sdram_controller.py:533" *)
                            casez (\$299 )
                              /* src = "sdram_controller.py:533" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$301 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$307 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                  (* src = "sdram_controller.py:613" *)
                                  casez (\$309 )
                                    /* src = "sdram_controller.py:613" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$311 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$313 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$315 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$317 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:352" *)
                                  casez (\$319 )
                                    /* src = "sdram_controller.py:352" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$321 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$323 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$325 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$327 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                          begin
                            (* src = "sdram_controller.py:546" *)
                            casez (\$329 )
                              /* src = "sdram_controller.py:546" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                            (* src = "sdram_controller.py:549" *)
                            casez (\$331 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$333 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:533" *)
                      casez (\$335 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramClkEn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    cmdRemainingCyclesCounter = 2'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$337 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$339 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$341 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$343 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:371" *)
                      casez (\$345 )
                        /* src = "sdram_controller.py:371" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:374" *)
                      casez (\$347 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$349 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$351 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$353 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$355 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$357 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                          begin
                            (* src = "sdram_controller.py:486" *)
                            casez (\$359 )
                              /* src = "sdram_controller.py:486" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:489" *)
                            casez (\$361 )
                              /* src = "sdram_controller.py:489" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$363 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$365 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                          begin
                            (* src = "sdram_controller.py:546" *)
                            casez (\$367 )
                              /* src = "sdram_controller.py:546" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:549" *)
                            casez (\$369 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$371 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$373 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$375 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
        begin
          (* src = "sdram_controller.py:505" *)
          casez (\$377 )
            /* src = "sdram_controller.py:505" */
            1'h1:
                cmdRemainingCyclesCounter = 2'h1;
          endcase
          (* src = "sdram_controller.py:508" *)
          casez (\$379 )
            /* src = "sdram_controller.py:508" */
            1'h1:
                cmdRemainingCyclesCounter = 2'h0;
          endcase
        end
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$381 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$391 , \$389 , \$387  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  cmdRemainingCyclesCounter = 2'h1;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$393 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$395 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$397 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$399 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$403 , \$401  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$409 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:443" *)
                                  casez (\$411 )
                                    /* src = "sdram_controller.py:443" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$413 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$415 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$417 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$419 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$421 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$423 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$429 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:613" *)
                                  casez (\$431 )
                                    /* src = "sdram_controller.py:613" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:616" *)
                                  casez (\$433 )
                                    /* src = "sdram_controller.py:616" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$435 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                          begin
                            (* src = "sdram_controller.py:352" *)
                            casez (\$437 )
                              /* src = "sdram_controller.py:352" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:355" *)
                            casez (\$439 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$441 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$443 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$445 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$447 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$457 , \$455 , \$453  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  cmdRemainingCyclesCounter = 2'h1;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$459 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:505" *)
                      casez (\$461 )
                        /* src = "sdram_controller.py:505" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:508" *)
                      casez (\$463 )
                        /* src = "sdram_controller.py:508" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$465 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$467 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$473 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:399" *)
                                  casez (\$475 )
                                    /* src = "sdram_controller.py:399" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$477 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$479 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1020" *)
                      casez (\$481 )
                        /* src = "sdram_controller.py:1020" */
                        1'h1:
                          begin
                            (* src = "sdram_controller.py:533" *)
                            casez (\$483 )
                              /* src = "sdram_controller.py:533" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:536" *)
                            casez (\$485 )
                              /* src = "sdram_controller.py:536" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$487 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$493 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:613" *)
                                  casez (\$495 )
                                    /* src = "sdram_controller.py:613" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:616" *)
                                  casez (\$497 )
                                    /* src = "sdram_controller.py:616" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$499 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$501 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$503 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$505 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$507 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                begin
                                  (* src = "sdram_controller.py:352" *)
                                  casez (\$509 )
                                    /* src = "sdram_controller.py:352" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$511 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$513 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$515 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$517 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$519 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$521 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                          begin
                            (* src = "sdram_controller.py:546" *)
                            casez (\$523 )
                              /* src = "sdram_controller.py:546" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:549" *)
                            casez (\$525 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$527 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:533" *)
                      casez (\$529 )
                        /* src = "sdram_controller.py:533" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:536" *)
                      casez (\$531 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    cmdCompleted = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$533 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$535 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$537 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:386" *)
                      casez ({ \$541 , \$539  })
                        /* src = "sdram_controller.py:386" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:388" */
                        2'b1?:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$543 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$545 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$547 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$549 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                            (* src = "sdram_controller.py:497" *)
                            casez ({ \$553 , \$551  })
                              /* src = "sdram_controller.py:497" */
                              2'b?1:
                                  /* empty */;
                              /* src = "sdram_controller.py:499" */
                              2'b1?:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$555 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$557 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$559 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$561 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$563 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:508" *)
          casez (\$565 )
            /* src = "sdram_controller.py:508" */
            1'h1:
                cmdCompleted = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$567 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$577 , \$575 , \$573  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$579 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$581 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$583 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$587 , \$585  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$593 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$595 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$597 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$599 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$601 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$603 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$609 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                  (* src = "sdram_controller.py:616" *)
                                  casez (\$611 )
                                    /* src = "sdram_controller.py:616" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$613 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$615 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$617 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$619 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$621 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$631 , \$629 , \$627  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$633 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:508" *)
                      casez (\$635 )
                        /* src = "sdram_controller.py:508" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$637 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$639 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$645 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$647 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$649 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1020" *)
                      casez (\$651 )
                        /* src = "sdram_controller.py:1020" */
                        1'h1:
                            (* src = "sdram_controller.py:536" *)
                            casez (\$653 )
                              /* src = "sdram_controller.py:536" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$655 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$661 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                  (* src = "sdram_controller.py:616" *)
                                  casez (\$663 )
                                    /* src = "sdram_controller.py:616" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$665 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$667 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$669 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$671 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$673 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$675 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$677 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$679 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$681 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$683 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$685 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$687 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramCSn$next  = sdramCSn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$689 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$691 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$693 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$695 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \sdramCSn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$697 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$699 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$701 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$703 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                            (* src = "sdram_controller.py:489" *)
                            casez (\$705 )
                              /* src = "sdram_controller.py:489" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$707 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$709 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$711 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$713 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$715 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:508" *)
          casez (\$717 )
            /* src = "sdram_controller.py:508" */
            1'h1:
                \sdramCSn$next  = 1'h0;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$719 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$729 , \$727 , \$725  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$731 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$733 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$735 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$739 , \$737  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$745 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$747 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        \sdramCSn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$749 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$751 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$753 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$755 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$757 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$759 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$761 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$771 , \$769 , \$767  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$773 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:508" *)
                      casez (\$775 )
                        /* src = "sdram_controller.py:508" */
                        1'h1:
                            \sdramCSn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$777 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$779 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$785 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$787 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramCSn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$789 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* src = "sdram_controller.py:1020" *)
                      casez (\$791 )
                        /* src = "sdram_controller.py:1020" */
                        1'h1:
                            (* src = "sdram_controller.py:536" *)
                            casez (\$793 )
                              /* src = "sdram_controller.py:536" */
                              1'h1:
                                  \sdramCSn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$795 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$797 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$799 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$801 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$803 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        \sdramCSn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$805 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$807 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$809 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$811 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$813 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$815 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:536" *)
                      casez (\$817 )
                        /* src = "sdram_controller.py:536" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramCSn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    banksShouldRefresh = 1'h0;
    (* src = "sdram_controller.py:659" *)
    casez (bankController0_bankShouldRefresh)
      /* src = "sdram_controller.py:659" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
    (* src = "sdram_controller.py:659" *)
    casez (bankController1_bankShouldRefresh)
      /* src = "sdram_controller.py:659" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
    (* src = "sdram_controller.py:659" *)
    casez (bankController2_bankShouldRefresh)
      /* src = "sdram_controller.py:659" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
    (* src = "sdram_controller.py:659" *)
    casez (bankController3_bankShouldRefresh)
      /* src = "sdram_controller.py:659" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \repeatRefresh$next  = repeatRefresh;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$819 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \repeatRefresh$next  = 1'h0;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$821 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:739" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:739" */
                        1'h1:
                            \repeatRefresh$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:769" *)
                casez (\$823 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      (* src = "sdram_controller.py:772" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:772" */
                        1'h1:
                            \repeatRefresh$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \repeatRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \powerUpCounter$next  = powerUpCounter;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
              begin
                (* src = "sdram_controller.py:712" *)
                casez (\$825 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \powerUpCounter$next  = 15'h5dc0;
                      endcase
                endcase
                (* src = "sdram_controller.py:722" *)
                casez (\$827 )
                  /* src = "sdram_controller.py:722" */
                  1'h1:
                      (* src = "sdram_controller.py:723" *)
                      casez (\$829 )
                        /* src = "sdram_controller.py:723" */
                        1'h1:
                            \powerUpCounter$next  = \$832 [14:0];
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \powerUpCounter$next  = 15'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \cmdIndex$next  = cmdIndex;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
              begin
                (* src = "sdram_controller.py:712" *)
                casez (\$834 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \cmdIndex$next  = 4'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:722" *)
                casez (\$836 )
                  /* src = "sdram_controller.py:722" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:723" *)
                      casez (\$838 )
                        /* src = "sdram_controller.py:723" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:725" */
                        default:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$840 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:739" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:739" */
                        1'h1:
                            \cmdIndex$next  = 4'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:742" *)
                casez (\$842 )
                  /* src = "sdram_controller.py:742" */
                  1'h1:
                      (* src = "sdram_controller.py:744" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:744" */
                        1'h1:
                            \cmdIndex$next  = 4'h2;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$844 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:751" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:751" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$846 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* src = "sdram_controller.py:756" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:756" */
                        1'h1:
                            \cmdIndex$next  = 4'h4;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$848 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:760" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:760" */
                        1'h1:
                            \cmdIndex$next  = 4'h5;
                      endcase
                endcase
                (* src = "sdram_controller.py:763" *)
                casez (\$850 )
                  /* src = "sdram_controller.py:763" */
                  1'h1:
                      (* src = "sdram_controller.py:764" *)
                      casez ({ \$854 , \$852  })
                        /* src = "sdram_controller.py:764" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:766" */
                        2'b1?:
                            \cmdIndex$next  = 4'h6;
                      endcase
                endcase
                (* src = "sdram_controller.py:769" *)
                casez (\$856 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:772" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:772" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                        /* src = "sdram_controller.py:775" */
                        default:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:814" *)
                casez (\$858 )
                  /* src = "sdram_controller.py:814" */
                  1'h1:
                      \cmdIndex$next  = 4'h1;
                endcase
                (* src = "sdram_controller.py:820" *)
                casez (\$860 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:828" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:828" */
                              1'h1:
                                  \cmdIndex$next  = 4'h2;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:831" *)
                casez (\$862 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      (* src = "sdram_controller.py:834" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:834" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$864 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$868 , \$866  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* src = "sdram_controller.py:846" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:846" */
                              1'h1:
                                  \cmdIndex$next  = 4'h4;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:849" *)
                casez (\$870 )
                  /* src = "sdram_controller.py:849" */
                  1'h1:
                      (* src = "sdram_controller.py:851" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:851" */
                        1'h1:
                            \cmdIndex$next  = 4'h5;
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$872 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      \cmdIndex$next  = 4'h6;
                endcase
                (* src = "sdram_controller.py:862" *)
                casez (\$874 )
                  /* src = "sdram_controller.py:862" */
                  1'h1:
                      \cmdIndex$next  = 4'h7;
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$876 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:910" *)
                      casez (\$878 )
                        /* src = "sdram_controller.py:910" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:912" */
                        default:
                            \cmdIndex$next  = 4'h8;
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$880 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:924" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:924" */
                              1'h1:
                                  \cmdIndex$next  = 4'h9;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$882 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      (* src = "sdram_controller.py:929" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:929" */
                        1'h1:
                            \cmdIndex$next  = 4'ha;
                      endcase
                endcase
                (* src = "sdram_controller.py:932" *)
                casez (\$884 )
                  /* src = "sdram_controller.py:932" */
                  1'h1:
                      (* src = "sdram_controller.py:936" *)
                      casez (\$886 )
                        /* src = "sdram_controller.py:936" */
                        1'h1:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:951" *)
                casez (\$888 )
                  /* src = "sdram_controller.py:951" */
                  1'h1:
                      \cmdIndex$next  = 4'h1;
                endcase
                (* src = "sdram_controller.py:955" *)
                casez (\$890 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:962" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:962" */
                              1'h1:
                                  \cmdIndex$next  = 4'h2;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$892 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:967" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:967" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$894 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$896 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* src = "sdram_controller.py:1011" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1011" */
                              1'h1:
                                  \cmdIndex$next  = 4'h4;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$898 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$900 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* src = "sdram_controller.py:1057" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1057" */
                              1'h1:
                                  \cmdIndex$next  = 4'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$902 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      (* src = "sdram_controller.py:1067" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1067" */
                        1'h1:
                            \cmdIndex$next  = 4'h6;
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$904 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1076" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1076" */
                        1'h1:
                            \cmdIndex$next  = 4'h7;
                      endcase
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$906 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      (* src = "sdram_controller.py:1082" *)
                      casez (\$908 )
                        /* src = "sdram_controller.py:1082" */
                        1'h1:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \cmdIndex$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramRASn$next  = sdramRASn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$910 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \sdramRASn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$912 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$914 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \sdramRASn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$916 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$918 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                            (* src = "sdram_controller.py:489" *)
                            casez (\$920 )
                              /* src = "sdram_controller.py:489" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$922 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$924 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$926 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:508" *)
          casez (\$928 )
            /* src = "sdram_controller.py:508" */
            1'h1:
                \sdramRASn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$930 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$940 , \$938 , \$936  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$942 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$946 , \$944  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$952 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$954 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        \sdramRASn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$956 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$958 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$960 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$970 , \$968 , \$966  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$972 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:508" *)
                      casez (\$974 )
                        /* src = "sdram_controller.py:508" */
                        1'h1:
                            \sdramRASn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$976 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$978 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$984 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$986 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramRASn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$988 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$990 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$992 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        \sdramRASn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1094" *)
                casez (\$994 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$996 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$998 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramRASn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramCASn$next  = sdramCASn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$1000 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \sdramCASn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1002 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1004 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \sdramCASn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$1006 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$1008 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                            (* src = "sdram_controller.py:489" *)
                            casez (\$1010 )
                              /* src = "sdram_controller.py:489" */
                              1'h1:
                                  \sdramCASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1012 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1014 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1016 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramCASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:508" *)
          casez (\$1018 )
            /* src = "sdram_controller.py:508" */
            1'h1:
                \sdramCASn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1020 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1030 , \$1028 , \$1026  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramCASn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$1032 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$1036 , \$1034  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$1042 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$1044 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        \sdramCASn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1046 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1048 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  \sdramCASn$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1050 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1060 , \$1058 , \$1056  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramCASn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$1062 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:508" *)
                      casez (\$1064 )
                        /* src = "sdram_controller.py:508" */
                        1'h1:
                            \sdramCASn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$1066 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$1068 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$1074 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$1076 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramCASn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1078 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1080 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1082 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        \sdramCASn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1094" *)
                casez (\$1084 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1086 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1088 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramCASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramCASn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramWEn$next  = sdramWEn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:712" *)
                casez (\$1090 )
                  /* src = "sdram_controller.py:712" */
                  1'h1:
                      (* src = "sdram_controller.py:714" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:714" */
                        1'h1:
                            \sdramWEn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1092 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1094 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \sdramWEn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$1096 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$1098 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                            (* src = "sdram_controller.py:489" *)
                            casez (\$1100 )
                              /* src = "sdram_controller.py:489" */
                              1'h1:
                                  \sdramWEn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1102 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1104 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1106 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:508" *)
          casez (\$1108 )
            /* src = "sdram_controller.py:508" */
            1'h1:
                \sdramWEn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1110 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1120 , \$1118 , \$1116  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$1122 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$1126 , \$1124  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$1132 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$1134 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        \sdramWEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1136 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1138 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  \sdramWEn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1140 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1150 , \$1148 , \$1146  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:965" *)
                casez (\$1152 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:508" *)
                      casez (\$1154 )
                        /* src = "sdram_controller.py:508" */
                        1'h1:
                            \sdramWEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$1156 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$1158 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$1164 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$1166 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramWEn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1168 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1170 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1172 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        \sdramWEn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1094" *)
                casez (\$1174 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1176 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1178 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramWEn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \delayCounter$next  = delayCounter;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:708" *)
          casez (errorState)
            /* src = "sdram_controller.py:708" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:711" */
            default:
                (* src = "sdram_controller.py:722" *)
                casez (\$1180 )
                  /* src = "sdram_controller.py:722" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:723" *)
                      casez (\$1182 )
                        /* src = "sdram_controller.py:723" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:725" */
                        default:
                            \delayCounter$next  = 4'hf;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1184 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1186 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \delayCounter$next  = 4'h1;
                      endcase
                      (* src = "sdram_controller.py:386" *)
                      casez ({ \$1190 , \$1188  })
                        /* src = "sdram_controller.py:386" */
                        2'b?1:
                            \delayCounter$next  = \$1193 [3:0];
                        /* src = "sdram_controller.py:388" */
                        2'b1?:
                            \delayCounter$next  = 4'hf;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$1195 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:483" *)
                      casez (\$1197 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:485" */
                        default:
                          begin
                            (* src = "sdram_controller.py:489" *)
                            casez (\$1199 )
                              /* src = "sdram_controller.py:489" */
                              1'h1:
                                  \delayCounter$next  = 4'h3;
                            endcase
                            (* src = "sdram_controller.py:497" *)
                            casez ({ \$1203 , \$1201  })
                              /* src = "sdram_controller.py:497" */
                              2'b?1:
                                  \delayCounter$next  = \$1206 [3:0];
                              /* src = "sdram_controller.py:499" */
                              2'b1?:
                                  \delayCounter$next  = 4'hf;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1208 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:760" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:760" */
                        1'h1:
                            \delayCounter$next  = 4'h6;
                      endcase
                endcase
                (* src = "sdram_controller.py:763" *)
                casez (\$1210 )
                  /* src = "sdram_controller.py:763" */
                  1'h1:
                      (* src = "sdram_controller.py:764" *)
                      casez ({ \$1214 , \$1212  })
                        /* src = "sdram_controller.py:764" */
                        2'b?1:
                            \delayCounter$next  = \$1217 [3:0];
                        /* src = "sdram_controller.py:766" */
                        2'b1?:
                            \delayCounter$next  = 4'hf;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:831" *)
                casez (\$1219 )
                  /* src = "sdram_controller.py:831" */
                  1'h1:
                      (* src = "sdram_controller.py:834" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:834" */
                        1'h1:
                            \delayCounter$next  = 4'h5;
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$1221 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$1225 , \$1223  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            \delayCounter$next  = \$1228 [3:0];
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            \delayCounter$next  = 4'hf;
                      endcase
                endcase
                (* src = "sdram_controller.py:926" *)
                casez (\$1230 )
                  /* src = "sdram_controller.py:926" */
                  1'h1:
                      (* src = "sdram_controller.py:929" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:929" */
                        1'h1:
                            \delayCounter$next  = 4'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:932" *)
                casez (\$1232 )
                  /* src = "sdram_controller.py:932" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:934" *)
                      casez (\$1234 )
                        /* src = "sdram_controller.py:934" */
                        1'h1:
                            \delayCounter$next  = \$1237 [3:0];
                      endcase
                      (* src = "sdram_controller.py:936" *)
                      casez (\$1239 )
                        /* src = "sdram_controller.py:936" */
                        1'h1:
                            \delayCounter$next  = 4'hf;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:965" *)
                casez (\$1241 )
                  /* src = "sdram_controller.py:965" */
                  1'h1:
                      (* src = "sdram_controller.py:967" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:967" */
                        1'h1:
                            \delayCounter$next  = 4'h5;
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$1243 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:997" *)
                      casez (\$1245 )
                        /* src = "sdram_controller.py:997" */
                        1'h1:
                            \delayCounter$next  = \$1248 [3:0];
                      endcase
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$1250 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            \delayCounter$next  = 4'hf;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$1252 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$1254 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* src = "sdram_controller.py:1057" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1057" */
                              1'h1:
                                  \delayCounter$next  = 4'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1063" *)
                casez (\$1256 )
                  /* src = "sdram_controller.py:1063" */
                  1'h1:
                      (* src = "sdram_controller.py:1065" *)
                      casez (\$1258 )
                        /* src = "sdram_controller.py:1065" */
                        1'h1:
                            \delayCounter$next  = \$1261 [3:0];
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1263 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1070" *)
                      casez (\$1265 )
                        /* src = "sdram_controller.py:1070" */
                        1'h1:
                            \delayCounter$next  = \$1268 [3:0];
                      endcase
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1270 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  \delayCounter$next  = 4'h1;
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1078" *)
                casez (\$1272 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1080" *)
                      casez (\$1274 )
                        /* src = "sdram_controller.py:1080" */
                        1'h1:
                            \delayCounter$next  = \$1277 [3:0];
                      endcase
                      (* src = "sdram_controller.py:1082" *)
                      casez (\$1279 )
                        /* src = "sdram_controller.py:1082" */
                        1'h1:
                            \delayCounter$next  = 4'hf;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$1281 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* src = "sdram_controller.py:1096" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1096" */
                        1'h1:
                            \delayCounter$next  = 4'h6;
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$1283 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$1289 , \$1285  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            \delayCounter$next  = \$1292 [3:0];
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \delayCounter$next  = 4'hf;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \delayCounter$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramAddress$next  = sdramAddress;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1294 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1296 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \sdramAddress$next [10] = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$1298 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:748" *)
                      casez (\$1300 )
                        /* src = "sdram_controller.py:748" */
                        1'h1:
                          begin
                            \sdramAddress$next [10] = 1'h0;
                            \sdramAddress$next [9] = 1'h0;
                            \sdramAddress$next [8:7] = 2'h0;
                            \sdramAddress$next [6:4] = 3'h3;
                            \sdramAddress$next [3] = 1'h0;
                            \sdramAddress$next [2:0] = 3'h7;
                          end
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1302 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1312 , \$1310 , \$1308  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramAddress$next  = targetRowAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$1314 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$1318 , \$1316  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$1324 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$1326 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        \sdramAddress$next  = { 3'h0, targetColumnAddress };
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1328 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1330 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  \sdramAddress$next [10] = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1332 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1342 , \$1340 , \$1338  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramAddress$next  = targetRowAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$1344 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$1346 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$1352 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$1354 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramAddress$next  = { 3'h0, targetColumnAddress };
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1356 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1358 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1360 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        \sdramAddress$next [10] = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramAddress$next  = 11'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController0_bankState$next  = bankController0_bankState;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1362 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1364 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \bankController0_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1366 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1368 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1370 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController0_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:769" *)
                casez (\$1372 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      \bankController0_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1374 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1384 , \$1382 , \$1380  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1386 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController0_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController0_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1388 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1390 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1392 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \bankController0_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1394 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1404 , \$1402 , \$1400  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1406 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController0_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController0_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1408 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1410 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1412 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        (* src = "sdram_controller.py:359" *)
                                        casez (\$1414 )
                                          /* src = "sdram_controller.py:359" */
                                          1'h1:
                                              \bankController0_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$1416 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1418 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1420 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController0_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$1422 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$1428 , \$1424  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \bankController0_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController0_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController1_bankState$next  = bankController1_bankState;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1430 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1432 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \bankController1_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1434 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1436 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1438 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController1_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:769" *)
                casez (\$1440 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      \bankController1_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1442 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1452 , \$1450 , \$1448  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1454 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController1_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController1_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1456 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1458 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1460 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \bankController1_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1462 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1472 , \$1470 , \$1468  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1474 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController1_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController1_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1476 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1478 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1480 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        (* src = "sdram_controller.py:359" *)
                                        casez (\$1482 )
                                          /* src = "sdram_controller.py:359" */
                                          1'h1:
                                              \bankController1_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$1484 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1486 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1488 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController1_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$1490 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$1496 , \$1492  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \bankController1_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController1_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:663" *)
    casez (targetBankAddress)
      2'h0:
          targetBankState = bankController0_bankState;
      2'h1:
          targetBankState = bankController1_bankState;
      2'h2:
          targetBankState = bankController2_bankState;
      2'h?:
          targetBankState = bankController3_bankState;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController2_bankState$next  = bankController2_bankState;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1498 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1500 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \bankController2_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1502 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1504 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1506 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController2_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:769" *)
                casez (\$1508 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      \bankController2_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1510 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1520 , \$1518 , \$1516  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1522 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController2_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController2_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1524 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1526 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1528 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \bankController2_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1530 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1540 , \$1538 , \$1536  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1542 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController2_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController2_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1544 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1546 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1548 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        (* src = "sdram_controller.py:359" *)
                                        casez (\$1550 )
                                          /* src = "sdram_controller.py:359" */
                                          1'h1:
                                              \bankController2_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$1552 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1554 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1556 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController2_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$1558 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$1564 , \$1560  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \bankController2_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController2_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController3_bankState$next  = bankController3_bankState;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:737" *)
                casez (\$1566 )
                  /* src = "sdram_controller.py:737" */
                  1'h1:
                      (* src = "sdram_controller.py:374" *)
                      casez (\$1568 )
                        /* src = "sdram_controller.py:374" */
                        1'h1:
                            \bankController3_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1570 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1572 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1574 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController3_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:769" *)
                casez (\$1576 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      \bankController3_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1578 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1588 , \$1586 , \$1584  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1590 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController3_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController3_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$1592 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      (* src = "sdram_controller.py:922" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:922" */
                        1'h1:
                            (* src = "sdram_controller.py:355" *)
                            casez (\$1594 )
                              /* src = "sdram_controller.py:355" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1596 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \bankController3_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1598 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1608 , \$1606 , \$1604  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1610 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:336" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:336" */
                                          1'h1:
                                              \bankController3_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:338" */
                                          default:
                                              \bankController3_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1069" *)
                casez (\$1612 )
                  /* src = "sdram_controller.py:1069" */
                  1'h1:
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1614 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            (* src = "sdram_controller.py:1073" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1073" */
                              1'h1:
                                  (* src = "sdram_controller.py:355" *)
                                  casez (\$1616 )
                                    /* src = "sdram_controller.py:355" */
                                    1'h1:
                                        (* src = "sdram_controller.py:359" *)
                                        casez (\$1618 )
                                          /* src = "sdram_controller.py:359" */
                                          1'h1:
                                              \bankController3_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$1620 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1622 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:545" */
                        default:
                            (* src = "sdram_controller.py:549" *)
                            casez (\$1624 )
                              /* src = "sdram_controller.py:549" */
                              1'h1:
                                  \bankController3_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$1626 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$1632 , \$1628  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \bankController3_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController3_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \errorState$next  = errorState;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
              begin
                (* src = "sdram_controller.py:746" *)
                casez (\$1634 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:483" *)
                      casez (\$1636 )
                        /* src = "sdram_controller.py:483" */
                        1'h1:
                            \errorState$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:754" *)
                casez (\$1638 )
                  /* src = "sdram_controller.py:754" */
                  1'h1:
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1640 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            \errorState$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1642 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1652 , \$1650 , \$1648  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$1654 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$1658 , \$1656  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* src = "sdram_controller.py:439" *)
                            casez (\$1664 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$1666 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$1668 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            (* src = "sdram_controller.py:609" *)
                            casez (\$1674 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1676 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1686 , \$1684 , \$1682  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$1688 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$1690 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* src = "sdram_controller.py:395" *)
                            casez (\$1696 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$1698 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$1700 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* src = "sdram_controller.py:609" *)
                            casez (\$1706 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1094" *)
                casez (\$1708 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* src = "sdram_controller.py:543" *)
                      casez (\$1710 )
                        /* src = "sdram_controller.py:543" */
                        1'h1:
                            \errorState$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \errorState$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramBank$next  = sdramBank;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
                (* src = "sdram_controller.py:746" *)
                casez (\$1712 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:748" *)
                      casez (\$1714 )
                        /* src = "sdram_controller.py:748" */
                        1'h1:
                            \sdramBank$next  = 2'h0;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$1716 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1726 , \$1724 , \$1722  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramBank$next  = targetBankAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:837" *)
                casez (\$1728 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$1732 , \$1730  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:439" *)
                            casez (\$1738 )
                              /* src = "sdram_controller.py:439" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:442" */
                              default:
                                  (* src = "sdram_controller.py:446" *)
                                  casez (\$1740 )
                                    /* src = "sdram_controller.py:446" */
                                    1'h1:
                                        \sdramBank$next  = targetBankAddress;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$1742 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1752 , \$1750 , \$1748  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  \sdramBank$next  = targetBankAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$1754 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$1756 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$1762 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$1764 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramBank$next  = targetBankAddress;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramBank$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \burstWritesMode$next  = burstWritesMode;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
                (* src = "sdram_controller.py:746" *)
                casez (\$1766 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:751" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:751" */
                        1'h1:
                            \burstWritesMode$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \burstWritesMode$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlReady$next  = ctrlReady;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:733" *)
          casez (errorState)
            /* src = "sdram_controller.py:733" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:736" */
            default:
                (* src = "sdram_controller.py:769" *)
                casez (\$1768 )
                  /* src = "sdram_controller.py:769" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:772" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:772" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:775" */
                        default:
                            \ctrlReady$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:784" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:784" */
            2'b?1:
                /* empty */;
            /* src = "sdram_controller.py:787" */
            2'b1?:
                (* src = "sdram_controller.py:788" *)
                casez ({ \$1770 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:788" */
                  3'b??1:
                      /* empty */;
                  /* src = "sdram_controller.py:791" */
                  3'b?1?:
                      \ctrlReady$next  = 1'h0;
                  /* src = "sdram_controller.py:797" */
                  3'b1??:
                      \ctrlReady$next  = 1'h0;
                endcase
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:932" *)
                casez (\$1772 )
                  /* src = "sdram_controller.py:932" */
                  1'h1:
                      (* src = "sdram_controller.py:936" *)
                      casez (\$1774 )
                        /* src = "sdram_controller.py:936" */
                        1'h1:
                            \ctrlReady$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:1078" *)
                casez (\$1776 )
                  /* src = "sdram_controller.py:1078" */
                  1'h1:
                      (* src = "sdram_controller.py:1082" *)
                      casez (\$1778 )
                        /* src = "sdram_controller.py:1082" */
                        1'h1:
                            \ctrlReady$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlReady$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlAddress$next  = ctrlAddress;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          (* src = "sdram_controller.py:784" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:784" */
            2'b?1:
                /* empty */;
            /* src = "sdram_controller.py:787" */
            2'b1?:
                (* src = "sdram_controller.py:788" *)
                casez ({ \$1780 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:788" */
                  3'b??1:
                      /* empty */;
                  /* src = "sdram_controller.py:791" */
                  3'b?1?:
                      \ctrlAddress$next  = ctrlRdAddress;
                  /* src = "sdram_controller.py:797" */
                  3'b1??:
                      \ctrlAddress$next  = ctrlWrAddress;
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlAddress$next  = 21'h000000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \refreshRequired$next  = refreshRequired;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:814" *)
                casez (\$1782 )
                  /* src = "sdram_controller.py:814" */
                  1'h1:
                      \refreshRequired$next  = \$1792 ;
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:951" *)
                casez (\$1794 )
                  /* src = "sdram_controller.py:951" */
                  1'h1:
                      \refreshRequired$next  = \$1804 ;
                endcase
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
                (* src = "sdram_controller.py:1099" *)
                casez (\$1806 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$1812 , \$1808  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \refreshRequired$next  = 1'h0;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \refreshRequired$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController0_bankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1814 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1824 , \$1822 , \$1820  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1826 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController0_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1828 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1838 , \$1836 , \$1834  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1840 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController0_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController0_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1842 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1852 , \$1850 , \$1848  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1854 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController0_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1856 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1866 , \$1864 , \$1862  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1868 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController0_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:664" *)
    casez (targetBankAddress)
      2'h0:
          \targetBankCanActivate$next  = bankController0_bankCanActivate;
      2'h1:
          \targetBankCanActivate$next  = bankController1_bankCanActivate;
      2'h2:
          \targetBankCanActivate$next  = bankController2_bankCanActivate;
      2'h?:
          \targetBankCanActivate$next  = bankController3_bankCanActivate;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \targetBankCanActivate$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController1_bankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1870 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1880 , \$1878 , \$1876  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1882 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController1_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1884 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1894 , \$1892 , \$1890  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1896 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController1_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController1_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1898 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1908 , \$1906 , \$1904  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1910 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController1_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1912 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1922 , \$1920 , \$1918  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1924 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController1_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController2_bankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1926 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1936 , \$1934 , \$1932  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1938 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController2_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1940 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1950 , \$1948 , \$1946  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1952 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController2_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController2_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1954 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1964 , \$1962 , \$1960  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1966 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController2_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1968 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1978 , \$1976 , \$1974  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1980 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController2_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController3_bankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$1982 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$1992 , \$1990 , \$1988  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$1994 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController3_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$1996 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$2006 , \$2004 , \$2002  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$2008 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        bankController3_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController3_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
                (* src = "sdram_controller.py:820" *)
                casez (\$2010 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$2020 , \$2018 , \$2016  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$2022 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController3_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
                (* src = "sdram_controller.py:955" *)
                casez (\$2024 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:325" *)
                            casez ({ \$2034 , \$2032 , \$2030  })
                              /* src = "sdram_controller.py:325" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:327" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:330" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:334" *)
                                  casez (\$2036 )
                                    /* src = "sdram_controller.py:334" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:340" */
                                    default:
                                        bankController3_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramDataMasks$next  = sdramDataMasks;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:820" *)
                casez (\$2038 )
                  /* src = "sdram_controller.py:820" */
                  1'h1:
                      (* src = "sdram_controller.py:822" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:822" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:826" */
                        2'b1?:
                            (* src = "sdram_controller.py:828" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:828" */
                              1'h1:
                                  \sdramDataMasks$next  = targetMask;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$2040 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* src = "sdram_controller.py:915" *)
                      casez (\$2042 )
                        /* src = "sdram_controller.py:915" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$2048 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                  (* src = "sdram_controller.py:616" *)
                                  casez (\$2050 )
                                    /* src = "sdram_controller.py:616" */
                                    1'h1:
                                        \sdramDataMasks$next  = 4'hf;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:955" *)
                casez (\$2052 )
                  /* src = "sdram_controller.py:955" */
                  1'h1:
                      (* src = "sdram_controller.py:956" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:956" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:960" */
                        2'b1?:
                            (* src = "sdram_controller.py:962" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:962" */
                              1'h1:
                                  \sdramDataMasks$next  = targetMask;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:970" *)
                casez (\$2054 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$2056 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:395" *)
                            casez (\$2062 )
                              /* src = "sdram_controller.py:395" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:398" */
                              default:
                                  (* src = "sdram_controller.py:402" *)
                                  casez (\$2064 )
                                    /* src = "sdram_controller.py:402" */
                                    1'h1:
                                        \sdramDataMasks$next  = targetMask;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$2066 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$2068 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:609" *)
                            casez (\$2074 )
                              /* src = "sdram_controller.py:609" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:612" */
                              default:
                                  (* src = "sdram_controller.py:616" *)
                                  casez (\$2076 )
                                    /* src = "sdram_controller.py:616" */
                                    1'h1:
                                        \sdramDataMasks$next  = 4'hf;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramDataMasks$next  = 4'hf;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \pageColumnIndex$next  = pageColumnIndex;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:837" *)
                casez (\$2078 )
                  /* src = "sdram_controller.py:837" */
                  1'h1:
                      (* src = "sdram_controller.py:838" *)
                      casez ({ \$2082 , \$2080  })
                        /* src = "sdram_controller.py:838" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:840" */
                        2'b1?:
                            (* src = "sdram_controller.py:846" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:846" */
                              1'h1:
                                  \pageColumnIndex$next  = targetColumnAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:869" *)
                casez (\$2084 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:910" *)
                      casez (\$2086 )
                        /* src = "sdram_controller.py:910" */
                        1'h1:
                            \pageColumnIndex$next  = \$2089 [7:0];
                        /* src = "sdram_controller.py:912" */
                        default:
                            \pageColumnIndex$next  = 8'h00;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:970" *)
                casez (\$2091 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$2093 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            \pageColumnIndex$next  = targetColumnAddress;
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$2095 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$2097 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            \pageColumnIndex$next  = \$2100 [7:0];
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \pageColumnIndex$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlRdInProgress$next  = ctrlRdInProgress;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:862" *)
                casez (\$2102 )
                  /* src = "sdram_controller.py:862" */
                  1'h1:
                      \ctrlRdInProgress$next  = 1'h1;
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$2104 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      \ctrlRdInProgress$next  = 1'h0;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlRdInProgress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlRdIncAddress$next  = ctrlRdIncAddress;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:869" *)
                casez (\$2106 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      \ctrlRdIncAddress$next  = 1'h1;
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$2108 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      \ctrlRdIncAddress$next  = 1'h0;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlRdIncAddress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:665" *)
    casez (targetBankAddress)
      2'h0:
          \targetBankCanPreCharge$next  = bankController0_bankCanPreCharge;
      2'h1:
          \targetBankCanPreCharge$next  = bankController1_bankCanPreCharge;
      2'h2:
          \targetBankCanPreCharge$next  = bankController2_bankCanPreCharge;
      2'h?:
          \targetBankCanPreCharge$next  = bankController3_bankCanPreCharge;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \targetBankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    ctrlRdDataOut = 24'h000000;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:810" *)
          casez (errorState)
            /* src = "sdram_controller.py:810" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:813" */
            default:
              begin
                (* src = "sdram_controller.py:869" *)
                casez (\$2110 )
                  /* src = "sdram_controller.py:869" */
                  1'h1:
                      ctrlRdDataOut = sdramDqOut[23:0];
                endcase
                (* src = "sdram_controller.py:917" *)
                casez (\$2112 )
                  /* src = "sdram_controller.py:917" */
                  1'h1:
                      ctrlRdDataOut = sdramDqOut[23:0];
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlWrIncAddress$next  = ctrlWrIncAddress;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:970" *)
                casez (\$2114 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:997" *)
                      casez (\$2116 )
                        /* src = "sdram_controller.py:997" */
                        1'h1:
                            (* src = "sdram_controller.py:999" *)
                            casez (\$2118 )
                              /* src = "sdram_controller.py:999" */
                              1'h1:
                                  \ctrlWrIncAddress$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$2120 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* src = "sdram_controller.py:1061" *)
                      casez (\$2122 )
                        /* src = "sdram_controller.py:1061" */
                        1'h1:
                            \ctrlWrIncAddress$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlWrIncAddress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramDqWRn$next  = sdramDqWRn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:970" *)
                casez (\$2124 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$2126 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            \sdramDqWRn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$2128 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$2130 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            \sdramDqWRn$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramDqWRn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramDqIn$next  = sdramDqIn;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:970" *)
                casez (\$2132 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$2134 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            \sdramDqIn$next [23:0] = ctrlWrDataIn;
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$2136 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      \sdramDqIn$next [23:0] = ctrlWrDataIn;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramDqIn$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlWrInProgress$next  = ctrlWrInProgress;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:947" *)
          casez (errorState)
            /* src = "sdram_controller.py:947" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:950" */
            default:
              begin
                (* src = "sdram_controller.py:970" *)
                casez (\$2138 )
                  /* src = "sdram_controller.py:970" */
                  1'h1:
                      (* src = "sdram_controller.py:1001" *)
                      casez (\$2140 )
                        /* src = "sdram_controller.py:1001" */
                        1'h1:
                            \ctrlWrInProgress$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1013" *)
                casez (\$2142 )
                  /* src = "sdram_controller.py:1013" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1052" *)
                      casez (\$2144 )
                        /* src = "sdram_controller.py:1052" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1054" */
                        default:
                            (* src = "sdram_controller.py:1057" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1057" */
                              1'h1:
                                  \ctrlWrInProgress$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlWrInProgress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \refreshCmdIndex$next  = refreshCmdIndex;
    (* src = "sdram_controller.py:704" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:705" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:730" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:780" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:805" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:941" */
      3'h6:
          /* empty */;
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1087" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1090" *)
          casez (errorState)
            /* src = "sdram_controller.py:1090" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1093" */
            default:
              begin
                (* src = "sdram_controller.py:1094" *)
                casez (\$2146 )
                  /* src = "sdram_controller.py:1094" */
                  1'h1:
                      (* src = "sdram_controller.py:1096" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1096" */
                        1'h1:
                            \refreshCmdIndex$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1099" *)
                casez (\$2148 )
                  /* src = "sdram_controller.py:1099" */
                  1'h1:
                      (* src = "sdram_controller.py:1101" *)
                      casez ({ \$2154 , \$2150  })
                        /* src = "sdram_controller.py:1101" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1103" */
                        2'b1?:
                            \refreshCmdIndex$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \refreshCmdIndex$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:666" *)
    casez (targetBankAddress)
      2'h0:
          \targetBankRefreshCounter$next  = bankController0_bankREFIcyclesCounter;
      2'h1:
          \targetBankRefreshCounter$next  = bankController1_bankREFIcyclesCounter;
      2'h2:
          \targetBankRefreshCounter$next  = bankController2_bankREFIcyclesCounter;
      2'h?:
          \targetBankRefreshCounter$next  = bankController3_bankREFIcyclesCounter;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \targetBankRefreshCounter$next  = 10'h000;
    endcase
  end
  assign \$831  = \$832 ;
  assign \$1192  = \$1193 ;
  assign \$1205  = \$1206 ;
  assign \$1216  = \$1217 ;
  assign \$1227  = \$1228 ;
  assign \$1236  = \$1237 ;
  assign \$1247  = \$1248 ;
  assign \$1260  = \$1261 ;
  assign \$1267  = \$1268 ;
  assign \$1276  = \$1277 ;
  assign \$1291  = \$1292 ;
  assign \$2088  = \$2089 ;
  assign \$2099  = \$2100 ;
  assign clkSDRAM_clk = 1'h0;
  assign clkSDRAM_rst = 1'h0;
  assign targetMask = 4'h8;
  assign targetRowAddress = ctrlAddress[20:10];
  assign targetBankAddress = ctrlAddress[9:8];
  assign targetColumnAddress = ctrlAddress[7:0];
  assign sdramClk = 1'h0;
  assign \$33  = refreshCmdIndex;
  assign \$57  = refreshCmdIndex;
  assign \$121  = refreshCmdIndex;
  assign \$179  = refreshCmdIndex;
  assign \$205  = sdramClkEn;
  assign \$223  = sdramClkEn;
  assign \$277  = sdramClkEn;
  assign \$331  = sdramClkEn;
  assign \$333  = refreshCmdIndex;
  assign \$341  = sdramClkEn;
  assign \$347  = sdramClkEn;
  assign \$353  = sdramClkEn;
  assign \$361  = sdramClkEn;
  assign \$369  = sdramClkEn;
  assign \$375  = sdramClkEn;
  assign \$379  = sdramClkEn;
  assign \$391  = sdramClkEn;
  assign \$397  = sdramClkEn;
  assign \$413  = sdramClkEn;
  assign \$419  = sdramClkEn;
  assign \$433  = sdramClkEn;
  assign \$439  = sdramClkEn;
  assign \$445  = sdramClkEn;
  assign \$457  = sdramClkEn;
  assign \$463  = sdramClkEn;
  assign \$477  = sdramClkEn;
  assign \$485  = sdramClkEn;
  assign \$497  = sdramClkEn;
  assign \$503  = sdramClkEn;
  assign \$511  = sdramClkEn;
  assign \$517  = sdramClkEn;
  assign \$525  = sdramClkEn;
  assign \$527  = refreshCmdIndex;
  assign \$531  = sdramClkEn;
  assign \$535  = sdramClkEn;
  assign \$545  = sdramClkEn;
  assign \$559  = sdramClkEn;
  assign \$563  = sdramClkEn;
  assign \$565  = sdramClkEn;
  assign \$577  = sdramClkEn;
  assign \$581  = sdramClkEn;
  assign \$595  = sdramClkEn;
  assign \$599  = sdramClkEn;
  assign \$611  = sdramClkEn;
  assign \$615  = sdramClkEn;
  assign \$619  = sdramClkEn;
  assign \$631  = sdramClkEn;
  assign \$635  = sdramClkEn;
  assign \$647  = sdramClkEn;
  assign \$653  = sdramClkEn;
  assign \$663  = sdramClkEn;
  assign \$667  = sdramClkEn;
  assign \$673  = sdramClkEn;
  assign \$677  = sdramClkEn;
  assign \$683  = sdramClkEn;
  assign \$685  = refreshCmdIndex;
  assign \$687  = sdramClkEn;
  assign \$691  = sdramClkEn;
  assign \$695  = sdramClkEn;
  assign \$699  = sdramClkEn;
  assign \$705  = sdramClkEn;
  assign \$711  = sdramClkEn;
  assign \$715  = sdramClkEn;
  assign \$717  = sdramClkEn;
  assign \$729  = sdramClkEn;
  assign \$733  = sdramClkEn;
  assign \$747  = sdramClkEn;
  assign \$751  = sdramClkEn;
  assign \$755  = sdramClkEn;
  assign \$759  = sdramClkEn;
  assign \$771  = sdramClkEn;
  assign \$775  = sdramClkEn;
  assign \$787  = sdramClkEn;
  assign \$793  = sdramClkEn;
  assign \$797  = sdramClkEn;
  assign \$803  = sdramClkEn;
  assign \$807  = sdramClkEn;
  assign \$813  = sdramClkEn;
  assign \$815  = refreshCmdIndex;
  assign \$817  = sdramClkEn;
  assign \$914  = sdramClkEn;
  assign \$920  = sdramClkEn;
  assign \$926  = sdramClkEn;
  assign \$928  = sdramClkEn;
  assign \$940  = sdramClkEn;
  assign \$954  = sdramClkEn;
  assign \$958  = sdramClkEn;
  assign \$970  = sdramClkEn;
  assign \$974  = sdramClkEn;
  assign \$986  = sdramClkEn;
  assign \$992  = sdramClkEn;
  assign \$998  = sdramClkEn;
  assign \$1004  = sdramClkEn;
  assign \$1010  = sdramClkEn;
  assign \$1016  = sdramClkEn;
  assign \$1018  = sdramClkEn;
  assign \$1030  = sdramClkEn;
  assign \$1044  = sdramClkEn;
  assign \$1048  = sdramClkEn;
  assign \$1060  = sdramClkEn;
  assign \$1064  = sdramClkEn;
  assign \$1076  = sdramClkEn;
  assign \$1082  = sdramClkEn;
  assign \$1088  = sdramClkEn;
  assign \$1094  = sdramClkEn;
  assign \$1100  = sdramClkEn;
  assign \$1106  = sdramClkEn;
  assign \$1108  = sdramClkEn;
  assign \$1120  = sdramClkEn;
  assign \$1134  = sdramClkEn;
  assign \$1138  = sdramClkEn;
  assign \$1150  = sdramClkEn;
  assign \$1154  = sdramClkEn;
  assign \$1166  = sdramClkEn;
  assign \$1172  = sdramClkEn;
  assign \$1178  = sdramClkEn;
  assign \$1186  = sdramClkEn;
  assign \$1199  = sdramClkEn;
  assign \$1283  = refreshCmdIndex;
  assign \$1296  = sdramClkEn;
  assign \$1312  = sdramClkEn;
  assign \$1326  = sdramClkEn;
  assign \$1330  = sdramClkEn;
  assign \$1342  = sdramClkEn;
  assign \$1354  = sdramClkEn;
  assign \$1360  = sdramClkEn;
  assign \$1364  = sdramClkEn;
  assign \$1370  = sdramClkEn;
  assign \$1384  = sdramClkEn;
  assign \$1390  = sdramClkEn;
  assign \$1404  = sdramClkEn;
  assign \$1412  = sdramClkEn;
  assign \$1420  = sdramClkEn;
  assign \$1422  = refreshCmdIndex;
  assign \$1432  = sdramClkEn;
  assign \$1438  = sdramClkEn;
  assign \$1452  = sdramClkEn;
  assign \$1458  = sdramClkEn;
  assign \$1472  = sdramClkEn;
  assign \$1480  = sdramClkEn;
  assign \$1488  = sdramClkEn;
  assign \$1490  = refreshCmdIndex;
  assign \$1500  = sdramClkEn;
  assign \$1506  = sdramClkEn;
  assign \$1520  = sdramClkEn;
  assign \$1526  = sdramClkEn;
  assign \$1540  = sdramClkEn;
  assign \$1548  = sdramClkEn;
  assign \$1556  = sdramClkEn;
  assign \$1558  = refreshCmdIndex;
  assign \$1568  = sdramClkEn;
  assign \$1574  = sdramClkEn;
  assign \$1588  = sdramClkEn;
  assign \$1594  = sdramClkEn;
  assign \$1608  = sdramClkEn;
  assign \$1616  = sdramClkEn;
  assign \$1624  = sdramClkEn;
  assign \$1626  = refreshCmdIndex;
  assign \$1652  = sdramClkEn;
  assign \$1686  = sdramClkEn;
  assign \$1726  = sdramClkEn;
  assign \$1740  = sdramClkEn;
  assign \$1752  = sdramClkEn;
  assign \$1764  = sdramClkEn;
  assign \$1786  = { 1'h0, \$1784  };
  assign \$1798  = { 1'h0, \$1796  };
  assign \$1806  = refreshCmdIndex;
  assign \$1824  = sdramClkEn;
  assign \$1838  = sdramClkEn;
  assign \$1852  = sdramClkEn;
  assign \$1866  = sdramClkEn;
  assign \$1880  = sdramClkEn;
  assign \$1894  = sdramClkEn;
  assign \$1908  = sdramClkEn;
  assign \$1922  = sdramClkEn;
  assign \$1936  = sdramClkEn;
  assign \$1950  = sdramClkEn;
  assign \$1964  = sdramClkEn;
  assign \$1978  = sdramClkEn;
  assign \$1992  = sdramClkEn;
  assign \$2006  = sdramClkEn;
  assign \$2020  = sdramClkEn;
  assign \$2034  = sdramClkEn;
  assign \$2050  = sdramClkEn;
  assign \$2064  = sdramClkEn;
  assign \$2076  = sdramClkEn;
  assign \$2148  = refreshCmdIndex;
endmodule

(* \amaranth.hierarchy  = "top" *)
(* top =  1  *)
(* generator = "Amaranth" *)
module top(sdramClkEn, sdramRASn, sdramCASn, sdramWEn, sdramCSn, sdramAddress, sdramBank, sdramDqOut, sdramDqIn, sdramDqWRn, sdramDataMasks, ctrlReady, ctrlWrAddress, ctrlWr, ctrlWrDataIn, ctrlWrIncAddress, ctrlRdAddress, ctrlRd, ctrlRdDataOut, ctrlRdIncAddress, sdramClk
);
  (* src = "sdram_controller.py:218" *)
  input ctrlRd;
  wire ctrlRd;
  (* src = "sdram_controller.py:217" *)
  input [20:0] ctrlRdAddress;
  wire [20:0] ctrlRdAddress;
  (* src = "sdram_controller.py:219" *)
  output [23:0] ctrlRdDataOut;
  wire [23:0] ctrlRdDataOut;
  (* src = "sdram_controller.py:220" *)
  output ctrlRdIncAddress;
  wire ctrlRdIncAddress;
  (* src = "sdram_controller.py:209" *)
  output ctrlReady;
  wire ctrlReady;
  (* src = "sdram_controller.py:212" *)
  input ctrlWr;
  wire ctrlWr;
  (* src = "sdram_controller.py:211" *)
  input [20:0] ctrlWrAddress;
  wire [20:0] ctrlWrAddress;
  (* src = "sdram_controller.py:213" *)
  input [23:0] ctrlWrDataIn;
  wire [23:0] ctrlWrDataIn;
  (* src = "sdram_controller.py:214" *)
  output ctrlWrIncAddress;
  wire ctrlWrIncAddress;
  (* src = "sdram_controller.py:201" *)
  output [10:0] sdramAddress;
  wire [10:0] sdramAddress;
  (* src = "sdram_controller.py:202" *)
  output [1:0] sdramBank;
  wire [1:0] sdramBank;
  (* src = "sdram_controller.py:198" *)
  output sdramCASn;
  wire sdramCASn;
  (* src = "sdram_controller.py:200" *)
  output sdramCSn;
  wire sdramCSn;
  (* src = "sdram_controller.py:195" *)
  output sdramClk;
  wire sdramClk;
  (* src = "sdram_controller.py:196" *)
  output sdramClkEn;
  wire sdramClkEn;
  (* src = "sdram_controller.py:206" *)
  output [3:0] sdramDataMasks;
  wire [3:0] sdramDataMasks;
  (* src = "sdram_controller.py:204" *)
  output [31:0] sdramDqIn;
  wire [31:0] sdramDqIn;
  (* src = "sdram_controller.py:203" *)
  input [31:0] sdramDqOut;
  wire [31:0] sdramDqOut;
  (* src = "sdram_controller.py:205" *)
  output sdramDqWRn;
  wire sdramDqWRn;
  (* src = "sdram_controller.py:197" *)
  output sdramRASn;
  wire sdramRASn;
  (* src = "sdram_controller.py:199" *)
  output sdramWEn;
  wire sdramWEn;
  sdramController sdramController (
    .ctrlRd(ctrlRd),
    .ctrlRdAddress(ctrlRdAddress),
    .ctrlRdDataOut(ctrlRdDataOut),
    .ctrlRdIncAddress(ctrlRdIncAddress),
    .ctrlReady(ctrlReady),
    .ctrlWr(ctrlWr),
    .ctrlWrAddress(ctrlWrAddress),
    .ctrlWrDataIn(ctrlWrDataIn),
    .ctrlWrIncAddress(ctrlWrIncAddress),
    .sdramAddress(sdramAddress),
    .sdramBank(sdramBank),
    .sdramCASn(sdramCASn),
    .sdramCSn(sdramCSn),
    .sdramClk(sdramClk),
    .sdramClkEn(sdramClkEn),
    .sdramDataMasks(sdramDataMasks),
    .sdramDqIn(sdramDqIn),
    .sdramDqOut(sdramDqOut),
    .sdramDqWRn(sdramDqWRn),
    .sdramRASn(sdramRASn),
    .sdramWEn(sdramWEn)
  );
endmodule

