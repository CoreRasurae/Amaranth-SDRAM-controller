// SPDX-License-Identifier: GPL-3.0-only
/*
 * EG4S20BG256 SDRAM controller
 *
 * Copyright (C) 2023 Luís Mendes <luis.p.mendes@gmail.com>
 */
/* PageWords= 256, Address width: 8 *)
/* Number of Read/Write suspend cycles/wait states    : 0 *)
/* Row cycle time (same bank)                   - RC  : 8 */
/* RAS to CAS delay (same bank)                 - RCD : 3 */
/* PreCharge to Refresh/Row activate (same bank)- RP  : 3 */
/* Row activate to row activate (diff. banks)   - RRD : 2 */
/* Row activate to pre-charge cycles (same bank)- RAS : 6 */
/* Write recovery time                          - WR  : 1 */
/* Mode register set cycle cycles               - MRD : 2 */
/* Average refresh interval cycles              - REFI: 936 */
/* Mask bit offset                                    : 0 */
/* Column address width                               : 8 */
/* Bank address width                                 : 2 */
/* Row address width                                  : 11 */
/* Generated by Yosys 0.17+9 (git sha1 98c7804b8, clang 10.0.0-4ubuntu1 -fPIC -Os) */

(* \amaranth.hierarchy  = "top.sdramController.bankController0" *)
(* generator = "Amaranth" *)
module bankController0(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$1  = 0;
  (* src = "sdram_controller.py:1191" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1194" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1214" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1219" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1179" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1178" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1177" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1171" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1171" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1176" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1180" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1174" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1191" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1192" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1193" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1191" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1191" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1194" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1200" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$36  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1200" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1203" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1210" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1210" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1210" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1214" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1215" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1219" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1191" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1220" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1194" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1194" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1201" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1204" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* src = "sdram_controller.py:1201" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1212" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1212" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h7;
      /* src = "sdram_controller.py:1214" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1217" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1217" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1219" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController.bankController1" *)
(* generator = "Amaranth" *)
module bankController1(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$2  = 0;
  (* src = "sdram_controller.py:1191" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1194" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1214" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1219" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1179" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1178" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1177" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1171" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1171" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1176" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1180" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1174" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1191" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1192" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1193" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1191" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1191" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1194" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1200" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$36  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1200" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1203" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1210" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1210" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1210" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1214" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1215" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1219" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1191" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1220" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1194" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1194" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1201" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1204" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* src = "sdram_controller.py:1201" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1212" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1212" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h7;
      /* src = "sdram_controller.py:1214" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$2 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1217" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1217" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1219" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController.bankController2" *)
(* generator = "Amaranth" *)
module bankController2(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$3  = 0;
  (* src = "sdram_controller.py:1191" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1194" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1214" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1219" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1179" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1178" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1177" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1171" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1171" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1176" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1180" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1174" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1191" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1192" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1193" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1191" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1191" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1194" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1200" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$36  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1200" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1203" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1210" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1210" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1210" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1214" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1215" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1219" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1191" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1220" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1194" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1194" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1201" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1204" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* src = "sdram_controller.py:1201" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1212" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1212" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h7;
      /* src = "sdram_controller.py:1214" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$3 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1217" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1217" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1219" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController.bankController3" *)
(* generator = "Amaranth" *)
module bankController3(bankState, bankShouldRefresh, bankCanActivate, bankCanPreCharge, bankREFIcyclesCounter, bankActivated, otherBankActivated, clkSDRAM_rst, clkSDRAM_clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$4  = 0;
  (* src = "sdram_controller.py:1191" *)
  wire \$1 ;
  (* src = "sdram_controller.py:1192" *)
  wire \$11 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$13 ;
  (* src = "sdram_controller.py:1193" *)
  wire [10:0] \$14 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$16 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$18 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$20 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$22 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$24 ;
  (* src = "sdram_controller.py:1194" *)
  wire \$26 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$28 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$30 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$32 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$34 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$36 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$38 ;
  (* src = "sdram_controller.py:1200" *)
  wire \$40 ;
  (* src = "sdram_controller.py:1201" *)
  wire \$42 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$44 ;
  (* src = "sdram_controller.py:1203" *)
  wire [3:0] \$45 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$47 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$49 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$5 ;
  (* src = "sdram_controller.py:1210" *)
  wire \$51 ;
  (* src = "sdram_controller.py:1214" *)
  wire \$53 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$55 ;
  (* src = "sdram_controller.py:1215" *)
  wire [3:0] \$56 ;
  (* src = "sdram_controller.py:1219" *)
  wire \$58 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$60 ;
  (* src = "sdram_controller.py:1220" *)
  wire [1:0] \$61 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$7 ;
  (* src = "sdram_controller.py:1191" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1179" *)
  input bankActivated;
  wire bankActivated;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] bankActivatedCounter = 3'h0;
  (* src = "sdram_controller.py:1173" *)
  reg [2:0] \bankActivatedCounter$next ;
  (* src = "sdram_controller.py:1178" *)
  output bankCanActivate;
  wire bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  output bankCanPreCharge;
  reg bankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:1177" *)
  reg \bankCanPreCharge$next ;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] bankRAScyclesCounter = 3'h0;
  (* src = "sdram_controller.py:1172" *)
  reg [2:0] \bankRAScyclesCounter$next ;
  (* src = "sdram_controller.py:1171" *)
  output [9:0] bankREFIcyclesCounter;
  reg [9:0] bankREFIcyclesCounter = 10'h000;
  (* src = "sdram_controller.py:1171" *)
  reg [9:0] \bankREFIcyclesCounter$next ;
  (* src = "sdram_controller.py:1176" *)
  output bankShouldRefresh;
  reg bankShouldRefresh = 1'h0;
  (* src = "sdram_controller.py:1176" *)
  reg \bankShouldRefresh$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  input [2:0] bankState;
  wire [2:0] bankState;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_clk;
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1290" *)
  input clkSDRAM_rst;
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:1180" *)
  input otherBankActivated;
  wire otherBankActivated;
  (* src = "sdram_controller.py:1174" *)
  reg otherBankActivatedCounter = 1'h0;
  (* src = "sdram_controller.py:1174" *)
  reg \otherBankActivatedCounter$next ;
  assign \$9  = \$5  | (* src = "sdram_controller.py:1191" *) \$7 ;
  assign \$11  = bankREFIcyclesCounter > (* src = "sdram_controller.py:1192" *) 1'h0;
  assign \$14  = bankREFIcyclesCounter - (* src = "sdram_controller.py:1193" *) 1'h1;
  assign \$16  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$18  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$1  = bankState == (* src = "sdram_controller.py:1191" *) 1'h1;
  assign \$20  = \$16  | (* src = "sdram_controller.py:1191" *) \$18 ;
  assign \$22  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  assign \$24  = \$20  | (* src = "sdram_controller.py:1191" *) \$22 ;
  assign \$26  = bankREFIcyclesCounter <= (* src = "sdram_controller.py:1194" *) 2'h3;
  assign \$28  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$30  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$32  = \$28  | (* src = "sdram_controller.py:1200" *) \$30 ;
  assign \$34  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$36  = bankState == (* src = "sdram_controller.py:1200" *) 2'h2;
  assign \$38  = bankState == (* src = "sdram_controller.py:1200" *) 2'h3;
  assign \$3  = bankState == (* src = "sdram_controller.py:1191" *) 2'h2;
  assign \$40  = \$36  | (* src = "sdram_controller.py:1200" *) \$38 ;
  assign \$42  = bankRAScyclesCounter < (* src = "sdram_controller.py:1201" *) 3'h5;
  assign \$45  = bankRAScyclesCounter + (* src = "sdram_controller.py:1203" *) 1'h1;
  assign \$47  = ! (* src = "sdram_controller.py:1210" *) bankActivatedCounter;
  assign \$49  = ~ (* src = "sdram_controller.py:1210" *) otherBankActivatedCounter;
  assign \$51  = \$47  & (* src = "sdram_controller.py:1210" *) \$49 ;
  assign \$53  = bankActivatedCounter > (* src = "sdram_controller.py:1214" *) 1'h0;
  assign \$56  = bankActivatedCounter - (* src = "sdram_controller.py:1215" *) 1'h1;
  assign \$58  = otherBankActivatedCounter > (* src = "sdram_controller.py:1219" *) 1'h0;
  assign \$5  = \$1  | (* src = "sdram_controller.py:1191" *) \$3 ;
  assign \$61  = otherBankActivatedCounter - (* src = "sdram_controller.py:1220" *) 1'h1;
  always @(posedge clkSDRAM_clk)
    bankREFIcyclesCounter <= \bankREFIcyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankShouldRefresh <= \bankShouldRefresh$next ;
  always @(posedge clkSDRAM_clk)
    bankCanPreCharge <= \bankCanPreCharge$next ;
  always @(posedge clkSDRAM_clk)
    bankRAScyclesCounter <= \bankRAScyclesCounter$next ;
  always @(posedge clkSDRAM_clk)
    bankActivatedCounter <= \bankActivatedCounter$next ;
  always @(posedge clkSDRAM_clk)
    otherBankActivatedCounter <= \otherBankActivatedCounter$next ;
  assign \$7  = bankState == (* src = "sdram_controller.py:1191" *) 2'h3;
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankREFIcyclesCounter$next  = bankREFIcyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$9 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1192" *)
          casez (\$11 )
            /* src = "sdram_controller.py:1192" */
            1'h1:
                \bankREFIcyclesCounter$next  = \$14 [9:0];
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankREFIcyclesCounter$next  = 10'h3a7;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankREFIcyclesCounter$next  = 10'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankShouldRefresh$next  = bankShouldRefresh;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1191" *)
    casez (\$24 )
      /* src = "sdram_controller.py:1191" */
      1'h1:
          (* src = "sdram_controller.py:1194" *)
          casez (\$26 )
            /* src = "sdram_controller.py:1194" */
            1'h1:
                \bankShouldRefresh$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1196" */
      default:
          \bankShouldRefresh$next  = 1'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankShouldRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$32 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1201" *)
          casez (\$34 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankCanPreCharge$next  = 1'h0;
            /* src = "sdram_controller.py:1204" */
            default:
                \bankCanPreCharge$next  = 1'h1;
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankCanPreCharge$next  = 1'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankRAScyclesCounter$next  = bankRAScyclesCounter;
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:1200" *)
    casez (\$40 )
      /* src = "sdram_controller.py:1200" */
      1'h1:
          (* src = "sdram_controller.py:1201" *)
          casez (\$42 )
            /* src = "sdram_controller.py:1201" */
            1'h1:
                \bankRAScyclesCounter$next  = \$45 [2:0];
          endcase
      /* src = "sdram_controller.py:1206" */
      default:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankRAScyclesCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \bankActivatedCounter$next  = bankActivatedCounter;
    (* src = "sdram_controller.py:1212" *)
    casez ({ \$53 , bankActivated })
      /* src = "sdram_controller.py:1212" */
      2'b?1:
          \bankActivatedCounter$next  = 3'h7;
      /* src = "sdram_controller.py:1214" */
      2'b1?:
          \bankActivatedCounter$next  = \$56 [2:0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankActivatedCounter$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$4 ) begin end
    \otherBankActivatedCounter$next  = otherBankActivatedCounter;
    (* src = "sdram_controller.py:1217" *)
    casez ({ \$58 , otherBankActivated })
      /* src = "sdram_controller.py:1217" */
      2'b?1:
          \otherBankActivatedCounter$next  = 1'h1;
      /* src = "sdram_controller.py:1219" */
      2'b1?:
          \otherBankActivatedCounter$next  = \$61 [0];
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \otherBankActivatedCounter$next  = 1'h0;
    endcase
  end
  assign \$13  = \$14 ;
  assign \$44  = \$45 ;
  assign \$55  = \$56 ;
  assign \$60  = \$61 ;
  assign bankCanActivate = \$51 ;
endmodule

(* \amaranth.hierarchy  = "top.sdramController" *)
(* generator = "Amaranth" *)
module sdramController(sdramClkEn, sdramCSn, sdramRASn, sdramCASn, sdramWEn, sdramAddress, sdramBank, ctrlReady, ctrlRd, ctrlWr, ctrlRdAddress, ctrlWrAddress, sdramDataMasks, ctrlRdIncAddress, ctrlRdDataOut, sdramDqOut, ctrlWrIncAddress, sdramDqWRn, sdramDqIn, ctrlWrDataIn, sdramClk
);
  reg \$auto$verilog_backend.cc:2083:dump_module$5  = 0;
  (* src = "sdram_controller.py:659" *)
  wire \$1 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1000 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1002 ;
  (* src = "sdram_controller.py:487" *)
  wire \$1004 ;
  (* src = "sdram_controller.py:493" *)
  wire \$1006 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1008 ;
  (* src = "sdram_controller.py:973" *)
  wire \$101 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1010 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1012 ;
  (* src = "sdram_controller.py:512" *)
  wire \$1014 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1016 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1018 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1020 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1022 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1024 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1026 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1028 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$103 ;
  (* src = "sdram_controller.py:841" *)
  wire \$1030 ;
  (* src = "sdram_controller.py:843" *)
  wire \$1032 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1034 ;
  (* src = "sdram_controller.py:444" *)
  wire \$1036 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1038 ;
  (* src = "sdram_controller.py:450" *)
  wire \$1040 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1042 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1044 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1046 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1048 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$105 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1050 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1052 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1054 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1056 ;
  (* src = "sdram_controller.py:973" *)
  wire \$1058 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$1060 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1062 ;
  (* src = "sdram_controller.py:400" *)
  wire \$1064 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1066 ;
  (* src = "sdram_controller.py:406" *)
  wire \$1068 ;
  (* src = "sdram_controller.py:1022" *)
  wire \$107 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1070 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1072 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1074 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1076 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1078 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1080 ;
  (* src = "sdram_controller.py:716" *)
  wire \$1082 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1084 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1086 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1088 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$109 ;
  (* src = "sdram_controller.py:487" *)
  wire \$1090 ;
  (* src = "sdram_controller.py:493" *)
  wire \$1092 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1094 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1096 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1098 ;
  (* src = "sdram_controller.py:727" *)
  wire \$11 ;
  (* src = "sdram_controller.py:512" *)
  wire \$1100 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1102 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1104 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1106 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1108 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$111 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1110 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1112 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1114 ;
  (* src = "sdram_controller.py:841" *)
  wire \$1116 ;
  (* src = "sdram_controller.py:843" *)
  wire \$1118 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1120 ;
  (* src = "sdram_controller.py:444" *)
  wire \$1122 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1124 ;
  (* src = "sdram_controller.py:450" *)
  wire \$1126 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1128 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$113 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1130 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1132 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1134 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1136 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1138 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1140 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1142 ;
  (* src = "sdram_controller.py:973" *)
  wire \$1144 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$1146 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1148 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$115 ;
  (* src = "sdram_controller.py:400" *)
  wire \$1150 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1152 ;
  (* src = "sdram_controller.py:406" *)
  wire \$1154 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1156 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1158 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1160 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1162 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1164 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1166 ;
  (* src = "sdram_controller.py:726" *)
  wire \$1168 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$117 ;
  (* src = "sdram_controller.py:727" *)
  wire \$1170 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1172 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1174 ;
  (* src = "sdram_controller.py:390" *)
  wire \$1176 ;
  (* src = "sdram_controller.py:392" *)
  wire \$1178 ;
  (* src = "sdram_controller.py:391" *)
  wire [5:0] \$1180 ;
  (* src = "sdram_controller.py:391" *)
  wire [5:0] \$1181 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1183 ;
  (* src = "sdram_controller.py:487" *)
  wire \$1185 ;
  (* src = "sdram_controller.py:493" *)
  wire \$1187 ;
  (* src = "sdram_controller.py:501" *)
  wire \$1189 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$119 ;
  (* src = "sdram_controller.py:503" *)
  wire \$1191 ;
  (* src = "sdram_controller.py:502" *)
  wire [5:0] \$1193 ;
  (* src = "sdram_controller.py:502" *)
  wire [5:0] \$1194 ;
  (* src = "sdram_controller.py:762" *)
  wire \$1196 ;
  (* src = "sdram_controller.py:767" *)
  wire \$1198 ;
  (* src = "sdram_controller.py:768" *)
  wire \$1200 ;
  (* src = "sdram_controller.py:770" *)
  wire \$1202 ;
  (* src = "sdram_controller.py:769" *)
  wire [5:0] \$1204 ;
  (* src = "sdram_controller.py:769" *)
  wire [5:0] \$1205 ;
  (* src = "sdram_controller.py:834" *)
  wire \$1207 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1209 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$121 ;
  (* src = "sdram_controller.py:841" *)
  wire \$1211 ;
  (* src = "sdram_controller.py:843" *)
  wire \$1213 ;
  (* src = "sdram_controller.py:842" *)
  wire [5:0] \$1215 ;
  (* src = "sdram_controller.py:842" *)
  wire [5:0] \$1216 ;
  (* src = "sdram_controller.py:929" *)
  wire \$1218 ;
  (* src = "sdram_controller.py:935" *)
  wire \$1220 ;
  (* src = "sdram_controller.py:937" *)
  wire \$1222 ;
  (* src = "sdram_controller.py:938" *)
  wire [5:0] \$1224 ;
  (* src = "sdram_controller.py:938" *)
  wire [5:0] \$1225 ;
  (* src = "sdram_controller.py:939" *)
  wire \$1227 ;
  (* src = "sdram_controller.py:967" *)
  wire \$1229 ;
  (* src = "sdram_controller.py:716" *)
  wire \$123 ;
  (* src = "sdram_controller.py:973" *)
  wire \$1231 ;
  (* src = "sdram_controller.py:1000" *)
  wire \$1233 ;
  (* src = "sdram_controller.py:1001" *)
  wire [5:0] \$1235 ;
  (* src = "sdram_controller.py:1001" *)
  wire [5:0] \$1236 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$1238 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$1240 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$1242 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$1244 ;
  (* src = "sdram_controller.py:1067" *)
  wire \$1246 ;
  (* src = "sdram_controller.py:1068" *)
  wire [5:0] \$1248 ;
  (* src = "sdram_controller.py:1068" *)
  wire [5:0] \$1249 ;
  (* src = "sdram_controller.py:741" *)
  wire \$125 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1251 ;
  (* src = "sdram_controller.py:1072" *)
  wire \$1253 ;
  (* src = "sdram_controller.py:1073" *)
  wire [5:0] \$1255 ;
  (* src = "sdram_controller.py:1073" *)
  wire [5:0] \$1256 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1258 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$1260 ;
  (* src = "sdram_controller.py:1082" *)
  wire \$1262 ;
  (* src = "sdram_controller.py:1083" *)
  wire [5:0] \$1264 ;
  (* src = "sdram_controller.py:1083" *)
  wire [5:0] \$1265 ;
  (* src = "sdram_controller.py:1084" *)
  wire \$1267 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1269 ;
  (* src = "sdram_controller.py:746" *)
  wire \$127 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1271 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1273 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1275 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1277 ;
  (* src = "sdram_controller.py:1104" *)
  wire [5:0] \$1279 ;
  (* src = "sdram_controller.py:1104" *)
  wire [5:0] \$1280 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1282 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1284 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1286 ;
  (* src = "sdram_controller.py:752" *)
  wire \$1288 ;
  (* src = "sdram_controller.py:750" *)
  wire \$129 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1290 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1292 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1294 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1296 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1298 ;
  (* src = "sdram_controller.py:773" *)
  wire \$13 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1300 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1302 ;
  (* src = "sdram_controller.py:841" *)
  wire \$1304 ;
  (* src = "sdram_controller.py:843" *)
  wire \$1306 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1308 ;
  (* src = "sdram_controller.py:758" *)
  wire \$131 ;
  (* src = "sdram_controller.py:444" *)
  wire \$1310 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1312 ;
  (* src = "sdram_controller.py:450" *)
  wire \$1314 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1316 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1318 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1320 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1322 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1324 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1326 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1328 ;
  (* src = "sdram_controller.py:762" *)
  wire \$133 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1330 ;
  (* src = "sdram_controller.py:973" *)
  wire \$1332 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$1334 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1336 ;
  (* src = "sdram_controller.py:400" *)
  wire \$1338 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1340 ;
  (* src = "sdram_controller.py:406" *)
  wire \$1342 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1344 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1346 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1348 ;
  (* src = "sdram_controller.py:824" *)
  wire \$135 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1350 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1352 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1354 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1356 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1358 ;
  (* src = "sdram_controller.py:773" *)
  wire \$1360 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1362 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1364 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1366 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1368 ;
  (* src = "sdram_controller.py:834" *)
  wire \$137 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1370 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1372 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1374 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1376 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1378 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1380 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1382 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1384 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1386 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1388 ;
  (* src = "sdram_controller.py:840" *)
  wire \$139 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1390 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1392 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1394 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1396 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1398 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1400 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1402 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1404 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1406 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1408 ;
  (* src = "sdram_controller.py:841" *)
  wire \$141 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1410 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1412 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1414 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1416 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1418 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1420 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1422 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1424 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1426 ;
  (* src = "sdram_controller.py:773" *)
  wire \$1428 ;
  (* src = "sdram_controller.py:843" *)
  wire \$143 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1430 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1432 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1434 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1436 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1438 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1440 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1442 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1444 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1446 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1448 ;
  (* src = "sdram_controller.py:853" *)
  wire \$145 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1450 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1452 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1454 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1456 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1458 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1460 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1462 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1464 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1466 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1468 ;
  (* src = "sdram_controller.py:872" *)
  wire \$147 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1470 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1472 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1474 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1476 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1478 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1480 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1482 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1484 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1486 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1488 ;
  (* src = "sdram_controller.py:918" *)
  wire \$149 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1490 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1492 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1494 ;
  (* src = "sdram_controller.py:773" *)
  wire \$1496 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1498 ;
  (* src = "sdram_controller.py:801" *)
  wire \$15 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1500 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1502 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1504 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1506 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1508 ;
  (* src = "sdram_controller.py:920" *)
  wire \$151 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1510 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1512 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1514 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1516 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1518 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1520 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1522 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1524 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1526 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1528 ;
  (* src = "sdram_controller.py:929" *)
  wire \$153 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1530 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1532 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1534 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1536 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1538 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1540 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1542 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1544 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1546 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1548 ;
  (* src = "sdram_controller.py:958" *)
  wire \$155 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1550 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1552 ;
  (* src = "sdram_controller.py:741" *)
  wire \$1554 ;
  (* src = "sdram_controller.py:378" *)
  wire \$1556 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1558 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1560 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1562 ;
  (* src = "sdram_controller.py:773" *)
  wire \$1564 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1566 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1568 ;
  (* src = "sdram_controller.py:967" *)
  wire \$157 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1570 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1572 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1574 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1576 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1578 ;
  (* src = "sdram_controller.py:920" *)
  wire \$1580 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1582 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1584 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1586 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1588 ;
  (* src = "sdram_controller.py:973" *)
  wire \$159 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1590 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1592 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1594 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1596 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1598 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$1600 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$1602 ;
  (* src = "sdram_controller.py:359" *)
  wire \$1604 ;
  (* src = "sdram_controller.py:363" *)
  wire \$1606 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1608 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$161 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1610 ;
  (* src = "sdram_controller.py:553" *)
  wire \$1612 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1614 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1616 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1618 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1620 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1622 ;
  (* src = "sdram_controller.py:487" *)
  wire \$1624 ;
  (* src = "sdram_controller.py:758" *)
  wire \$1626 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1628 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$163 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1630 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1632 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1634 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1636 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1638 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1640 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1642 ;
  (* src = "sdram_controller.py:841" *)
  wire \$1644 ;
  (* src = "sdram_controller.py:843" *)
  wire \$1646 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1648 ;
  (* src = "sdram_controller.py:1022" *)
  wire \$165 ;
  (* src = "sdram_controller.py:444" *)
  wire \$1650 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1652 ;
  (* src = "sdram_controller.py:872" *)
  wire \$1654 ;
  (* src = "sdram_controller.py:918" *)
  wire \$1656 ;
  (* src = "sdram_controller.py:613" *)
  wire \$1658 ;
  (* src = "sdram_controller.py:614" *)
  wire \$1660 ;
  (* src = "sdram_controller.py:613" *)
  wire \$1662 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1664 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1666 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1668 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$167 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1670 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1672 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1674 ;
  (* src = "sdram_controller.py:973" *)
  wire \$1676 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$1678 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1680 ;
  (* src = "sdram_controller.py:400" *)
  wire \$1682 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1684 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$1686 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$1688 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$169 ;
  (* src = "sdram_controller.py:613" *)
  wire \$1690 ;
  (* src = "sdram_controller.py:614" *)
  wire \$1692 ;
  (* src = "sdram_controller.py:613" *)
  wire \$1694 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$1696 ;
  (* src = "sdram_controller.py:547" *)
  wire \$1698 ;
  (* src = "sdram_controller.py:799" *)
  wire \$17 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1700 ;
  (* src = "sdram_controller.py:752" *)
  wire \$1702 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1704 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1706 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1708 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$171 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1710 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1712 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1714 ;
  (* src = "sdram_controller.py:840" *)
  wire \$1716 ;
  (* src = "sdram_controller.py:841" *)
  wire \$1718 ;
  (* src = "sdram_controller.py:843" *)
  wire \$1720 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1722 ;
  (* src = "sdram_controller.py:444" *)
  wire \$1724 ;
  (* src = "sdram_controller.py:443" *)
  wire \$1726 ;
  (* src = "sdram_controller.py:450" *)
  wire \$1728 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$173 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1730 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1732 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1734 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1736 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1738 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1740 ;
  (* src = "sdram_controller.py:973" *)
  wire \$1742 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$1744 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1746 ;
  (* src = "sdram_controller.py:400" *)
  wire \$1748 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$175 ;
  (* src = "sdram_controller.py:399" *)
  wire \$1750 ;
  (* src = "sdram_controller.py:406" *)
  wire \$1752 ;
  (* src = "sdram_controller.py:750" *)
  wire \$1754 ;
  (* src = "sdram_controller.py:773" *)
  wire \$1756 ;
  (* src = "sdram_controller.py:801" *)
  wire \$1758 ;
  (* src = "sdram_controller.py:935" *)
  wire \$1760 ;
  (* src = "sdram_controller.py:939" *)
  wire \$1762 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$1764 ;
  (* src = "sdram_controller.py:1084" *)
  wire \$1766 ;
  (* src = "sdram_controller.py:801" *)
  wire \$1768 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$177 ;
  (* src = "sdram_controller.py:818" *)
  wire \$1770 ;
  (* src = "sdram_controller.py:822" *)
  wire [9:0] \$1772 ;
  (* src = "sdram_controller.py:822" *)
  wire [10:0] \$1774 ;
  (* src = "sdram_controller.py:822" *)
  wire [11:0] \$1776 ;
  (* src = "sdram_controller.py:822" *)
  wire [12:0] \$1778 ;
  (* src = "sdram_controller.py:822" *)
  wire \$1780 ;
  (* src = "sdram_controller.py:954" *)
  wire \$1782 ;
  (* src = "sdram_controller.py:956" *)
  wire [9:0] \$1784 ;
  (* src = "sdram_controller.py:956" *)
  wire [10:0] \$1786 ;
  (* src = "sdram_controller.py:956" *)
  wire [11:0] \$1788 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$179 ;
  (* src = "sdram_controller.py:956" *)
  wire [12:0] \$1790 ;
  (* src = "sdram_controller.py:956" *)
  wire \$1792 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$1794 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$1796 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1798 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$1800 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1802 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1804 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1806 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1808 ;
  (* src = "sdram_controller.py:716" *)
  wire \$181 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1810 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1812 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1814 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1816 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1818 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1820 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1822 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1824 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1826 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1828 ;
  (* src = "sdram_controller.py:537" *)
  wire \$183 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1830 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1832 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1834 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1836 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1838 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1840 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1842 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1844 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1846 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1848 ;
  (* src = "sdram_controller.py:741" *)
  wire \$185 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1850 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1852 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1854 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1856 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1858 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1860 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1862 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1864 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1866 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1868 ;
  (* src = "sdram_controller.py:375" *)
  wire \$187 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1870 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1872 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1874 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1876 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1878 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1880 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1882 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1884 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1886 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1888 ;
  (* src = "sdram_controller.py:746" *)
  wire \$189 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1890 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1892 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1894 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1896 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1898 ;
  (* src = "sdram_controller.py:805" *)
  wire \$19 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1900 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1902 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1904 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1906 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1908 ;
  (* src = "sdram_controller.py:537" *)
  wire \$191 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1910 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1912 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1914 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1916 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1918 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1920 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1922 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1924 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1926 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1928 ;
  (* src = "sdram_controller.py:750" *)
  wire \$193 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1930 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1932 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1934 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1936 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1938 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1940 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1942 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1944 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1946 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1948 ;
  (* src = "sdram_controller.py:487" *)
  wire \$195 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1950 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1952 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1954 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1956 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1958 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1960 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1962 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1964 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1966 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1968 ;
  (* src = "sdram_controller.py:490" *)
  wire \$197 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1970 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1972 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1974 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1976 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1978 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1980 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1982 ;
  (* src = "sdram_controller.py:958" *)
  wire \$1984 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1986 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1988 ;
  (* src = "sdram_controller.py:758" *)
  wire \$199 ;
  (* src = "sdram_controller.py:329" *)
  wire \$1990 ;
  (* src = "sdram_controller.py:331" *)
  wire \$1992 ;
  (* src = "sdram_controller.py:334" *)
  wire \$1994 ;
  (* src = "sdram_controller.py:338" *)
  wire \$1996 ;
  (* src = "sdram_controller.py:824" *)
  wire \$1998 ;
  (* src = "sdram_controller.py:329" *)
  wire \$2000 ;
  (* src = "sdram_controller.py:329" *)
  wire \$2002 ;
  (* src = "sdram_controller.py:329" *)
  wire \$2004 ;
  (* src = "sdram_controller.py:331" *)
  wire \$2006 ;
  (* src = "sdram_controller.py:334" *)
  wire \$2008 ;
  (* src = "sdram_controller.py:547" *)
  wire \$201 ;
  (* src = "sdram_controller.py:338" *)
  wire \$2010 ;
  (* src = "sdram_controller.py:958" *)
  wire \$2012 ;
  (* src = "sdram_controller.py:329" *)
  wire \$2014 ;
  (* src = "sdram_controller.py:329" *)
  wire \$2016 ;
  (* src = "sdram_controller.py:329" *)
  wire \$2018 ;
  (* src = "sdram_controller.py:331" *)
  wire \$2020 ;
  (* src = "sdram_controller.py:334" *)
  wire \$2022 ;
  (* src = "sdram_controller.py:338" *)
  wire \$2024 ;
  (* src = "sdram_controller.py:840" *)
  wire \$2026 ;
  (* src = "sdram_controller.py:841" *)
  wire \$2028 ;
  (* src = "sdram_controller.py:550" *)
  wire \$203 ;
  (* src = "sdram_controller.py:843" *)
  wire \$2030 ;
  (* src = "sdram_controller.py:920" *)
  wire \$2032 ;
  (* src = "sdram_controller.py:840" *)
  wire \$2034 ;
  (* src = "sdram_controller.py:841" *)
  wire \$2036 ;
  (* src = "sdram_controller.py:843" *)
  wire \$2038 ;
  (* src = "sdram_controller.py:872" *)
  wire \$2040 ;
  (* src = "sdram_controller.py:918" *)
  wire \$2042 ;
  (* src = "sdram_controller.py:613" *)
  wire \$2044 ;
  (* src = "sdram_controller.py:614" *)
  wire \$2046 ;
  (* src = "sdram_controller.py:613" *)
  wire \$2048 ;
  (* src = "sdram_controller.py:553" *)
  wire \$205 ;
  (* src = "sdram_controller.py:620" *)
  wire \$2050 ;
  (* src = "sdram_controller.py:973" *)
  wire \$2052 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$2054 ;
  (* src = "sdram_controller.py:399" *)
  wire \$2056 ;
  (* src = "sdram_controller.py:400" *)
  wire \$2058 ;
  (* src = "sdram_controller.py:399" *)
  wire \$2060 ;
  (* src = "sdram_controller.py:406" *)
  wire \$2062 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$2064 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$2066 ;
  (* src = "sdram_controller.py:613" *)
  wire \$2068 ;
  (* src = "sdram_controller.py:762" *)
  wire \$207 ;
  (* src = "sdram_controller.py:614" *)
  wire \$2070 ;
  (* src = "sdram_controller.py:613" *)
  wire \$2072 ;
  (* src = "sdram_controller.py:620" *)
  wire \$2074 ;
  (* src = "sdram_controller.py:853" *)
  wire \$2076 ;
  (* src = "sdram_controller.py:872" *)
  wire \$2078 ;
  (* src = "sdram_controller.py:913" *)
  wire \$2080 ;
  (* src = "sdram_controller.py:914" *)
  wire [8:0] \$2082 ;
  (* src = "sdram_controller.py:914" *)
  wire [8:0] \$2083 ;
  (* src = "sdram_controller.py:973" *)
  wire \$2085 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$2087 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$2089 ;
  (* src = "sdram_controller.py:537" *)
  wire \$209 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$2091 ;
  (* src = "sdram_controller.py:1055" *)
  wire [8:0] \$2093 ;
  (* src = "sdram_controller.py:1055" *)
  wire [8:0] \$2094 ;
  (* src = "sdram_controller.py:872" *)
  wire \$2096 ;
  (* src = "sdram_controller.py:920" *)
  wire \$2098 ;
  (* src = "sdram_controller.py:824" *)
  wire \$21 ;
  (* src = "sdram_controller.py:872" *)
  wire \$2100 ;
  (* src = "sdram_controller.py:920" *)
  wire \$2102 ;
  (* src = "sdram_controller.py:967" *)
  wire \$2104 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$2106 ;
  (* src = "sdram_controller.py:1063" *)
  wire \$2108 ;
  (* src = "sdram_controller.py:509" *)
  wire \$211 ;
  (* src = "sdram_controller.py:973" *)
  wire \$2110 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$2112 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$2114 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$2116 ;
  (* src = "sdram_controller.py:973" *)
  wire \$2118 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$2120 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$2122 ;
  (* src = "sdram_controller.py:217" *)
  wire [31:0] \$2124 ;
  (* src = "sdram_controller.py:973" *)
  wire \$2126 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$2128 ;
  (* src = "sdram_controller.py:824" *)
  wire \$213 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$2130 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$2132 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$2134 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$2136 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$2138 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$2140 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$2142 ;
  (* src = "sdram_controller.py:329" *)
  wire \$215 ;
  (* src = "sdram_controller.py:329" *)
  wire \$217 ;
  (* src = "sdram_controller.py:329" *)
  wire \$219 ;
  (* src = "sdram_controller.py:331" *)
  wire \$221 ;
  (* src = "sdram_controller.py:334" *)
  wire \$223 ;
  (* src = "sdram_controller.py:834" *)
  wire \$225 ;
  (* src = "sdram_controller.py:537" *)
  wire \$227 ;
  (* src = "sdram_controller.py:840" *)
  wire \$229 ;
  (* src = "sdram_controller.py:935" *)
  wire \$23 ;
  (* src = "sdram_controller.py:841" *)
  wire \$231 ;
  (* src = "sdram_controller.py:843" *)
  wire \$233 ;
  (* src = "sdram_controller.py:443" *)
  wire \$235 ;
  (* src = "sdram_controller.py:444" *)
  wire \$237 ;
  (* src = "sdram_controller.py:443" *)
  wire \$239 ;
  (* src = "sdram_controller.py:447" *)
  wire \$241 ;
  (* src = "sdram_controller.py:853" *)
  wire \$243 ;
  (* src = "sdram_controller.py:537" *)
  wire \$245 ;
  (* src = "sdram_controller.py:872" *)
  wire \$247 ;
  (* src = "sdram_controller.py:918" *)
  wire \$249 ;
  (* src = "sdram_controller.py:939" *)
  wire \$25 ;
  (* src = "sdram_controller.py:613" *)
  wire \$251 ;
  (* src = "sdram_controller.py:614" *)
  wire \$253 ;
  (* src = "sdram_controller.py:613" *)
  wire \$255 ;
  (* src = "sdram_controller.py:617" *)
  wire \$257 ;
  (* src = "sdram_controller.py:920" *)
  wire \$259 ;
  (* src = "sdram_controller.py:356" *)
  wire \$261 ;
  (* src = "sdram_controller.py:929" *)
  wire \$263 ;
  (* src = "sdram_controller.py:537" *)
  wire \$265 ;
  (* src = "sdram_controller.py:958" *)
  wire \$267 ;
  (* src = "sdram_controller.py:329" *)
  wire \$269 ;
  (* src = "sdram_controller.py:958" *)
  wire \$27 ;
  (* src = "sdram_controller.py:329" *)
  wire \$271 ;
  (* src = "sdram_controller.py:329" *)
  wire \$273 ;
  (* src = "sdram_controller.py:331" *)
  wire \$275 ;
  (* src = "sdram_controller.py:334" *)
  wire \$277 ;
  (* src = "sdram_controller.py:967" *)
  wire \$279 ;
  (* src = "sdram_controller.py:537" *)
  wire \$281 ;
  (* src = "sdram_controller.py:973" *)
  wire \$283 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$285 ;
  (* src = "sdram_controller.py:399" *)
  wire \$287 ;
  (* src = "sdram_controller.py:400" *)
  wire \$289 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$29 ;
  (* src = "sdram_controller.py:399" *)
  wire \$291 ;
  (* src = "sdram_controller.py:403" *)
  wire \$293 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$295 ;
  (* src = "sdram_controller.py:1022" *)
  wire \$297 ;
  (* src = "sdram_controller.py:537" *)
  wire \$299 ;
  (* src = "sdram_controller.py:659" *)
  wire \$3 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$301 ;
  (* src = "sdram_controller.py:613" *)
  wire \$303 ;
  (* src = "sdram_controller.py:614" *)
  wire \$305 ;
  (* src = "sdram_controller.py:613" *)
  wire \$307 ;
  (* src = "sdram_controller.py:617" *)
  wire \$309 ;
  (* src = "sdram_controller.py:1084" *)
  wire \$31 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$311 ;
  (* src = "sdram_controller.py:537" *)
  wire \$313 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$315 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$317 ;
  (* src = "sdram_controller.py:356" *)
  wire \$319 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$321 ;
  (* src = "sdram_controller.py:537" *)
  wire \$323 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$325 ;
  (* src = "sdram_controller.py:547" *)
  wire \$327 ;
  (* src = "sdram_controller.py:550" *)
  wire \$329 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$33 ;
  (* src = "sdram_controller.py:553" *)
  wire \$331 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$333 ;
  (* src = "sdram_controller.py:537" *)
  wire \$335 ;
  (* src = "sdram_controller.py:716" *)
  wire \$337 ;
  (* src = "sdram_controller.py:537" *)
  wire \$339 ;
  (* src = "sdram_controller.py:540" *)
  wire \$341 ;
  (* src = "sdram_controller.py:741" *)
  wire \$343 ;
  (* src = "sdram_controller.py:375" *)
  wire \$345 ;
  (* src = "sdram_controller.py:378" *)
  wire \$347 ;
  (* src = "sdram_controller.py:746" *)
  wire \$349 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$35 ;
  (* src = "sdram_controller.py:537" *)
  wire \$351 ;
  (* src = "sdram_controller.py:540" *)
  wire \$353 ;
  (* src = "sdram_controller.py:750" *)
  wire \$355 ;
  (* src = "sdram_controller.py:487" *)
  wire \$357 ;
  (* src = "sdram_controller.py:490" *)
  wire \$359 ;
  (* src = "sdram_controller.py:493" *)
  wire \$361 ;
  (* src = "sdram_controller.py:758" *)
  wire \$363 ;
  (* src = "sdram_controller.py:547" *)
  wire \$365 ;
  (* src = "sdram_controller.py:550" *)
  wire \$367 ;
  (* src = "sdram_controller.py:553" *)
  wire \$369 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$37 ;
  (* src = "sdram_controller.py:762" *)
  wire \$371 ;
  (* src = "sdram_controller.py:537" *)
  wire \$373 ;
  (* src = "sdram_controller.py:540" *)
  wire \$375 ;
  (* src = "sdram_controller.py:509" *)
  wire \$377 ;
  (* src = "sdram_controller.py:512" *)
  wire \$379 ;
  (* src = "sdram_controller.py:824" *)
  wire \$381 ;
  (* src = "sdram_controller.py:329" *)
  wire \$383 ;
  (* src = "sdram_controller.py:329" *)
  wire \$385 ;
  (* src = "sdram_controller.py:329" *)
  wire \$387 ;
  (* src = "sdram_controller.py:331" *)
  wire \$389 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$39 ;
  (* src = "sdram_controller.py:334" *)
  wire \$391 ;
  (* src = "sdram_controller.py:834" *)
  wire \$393 ;
  (* src = "sdram_controller.py:537" *)
  wire \$395 ;
  (* src = "sdram_controller.py:540" *)
  wire \$397 ;
  (* src = "sdram_controller.py:840" *)
  wire \$399 ;
  (* src = "sdram_controller.py:841" *)
  wire \$401 ;
  (* src = "sdram_controller.py:843" *)
  wire \$403 ;
  (* src = "sdram_controller.py:443" *)
  wire \$405 ;
  (* src = "sdram_controller.py:444" *)
  wire \$407 ;
  (* src = "sdram_controller.py:443" *)
  wire \$409 ;
  (* src = "sdram_controller.py:1112" *)
  wire \$41 ;
  (* src = "sdram_controller.py:447" *)
  wire \$411 ;
  (* src = "sdram_controller.py:450" *)
  wire \$413 ;
  (* src = "sdram_controller.py:853" *)
  wire \$415 ;
  (* src = "sdram_controller.py:537" *)
  wire \$417 ;
  (* src = "sdram_controller.py:540" *)
  wire \$419 ;
  (* src = "sdram_controller.py:872" *)
  wire \$421 ;
  (* src = "sdram_controller.py:918" *)
  wire \$423 ;
  (* src = "sdram_controller.py:613" *)
  wire \$425 ;
  (* src = "sdram_controller.py:614" *)
  wire \$427 ;
  (* src = "sdram_controller.py:613" *)
  wire \$429 ;
  (* src = "sdram_controller.py:1114" *)
  wire \$43 ;
  (* src = "sdram_controller.py:617" *)
  wire \$431 ;
  (* src = "sdram_controller.py:620" *)
  wire \$433 ;
  (* src = "sdram_controller.py:920" *)
  wire \$435 ;
  (* src = "sdram_controller.py:356" *)
  wire \$437 ;
  (* src = "sdram_controller.py:359" *)
  wire \$439 ;
  (* src = "sdram_controller.py:929" *)
  wire \$441 ;
  (* src = "sdram_controller.py:537" *)
  wire \$443 ;
  (* src = "sdram_controller.py:540" *)
  wire \$445 ;
  (* src = "sdram_controller.py:958" *)
  wire \$447 ;
  (* src = "sdram_controller.py:329" *)
  wire \$449 ;
  (* src = "sdram_controller.py:726" *)
  wire \$45 ;
  (* src = "sdram_controller.py:329" *)
  wire \$451 ;
  (* src = "sdram_controller.py:329" *)
  wire \$453 ;
  (* src = "sdram_controller.py:331" *)
  wire \$455 ;
  (* src = "sdram_controller.py:334" *)
  wire \$457 ;
  (* src = "sdram_controller.py:967" *)
  wire \$459 ;
  (* src = "sdram_controller.py:537" *)
  wire \$461 ;
  (* src = "sdram_controller.py:540" *)
  wire \$463 ;
  (* src = "sdram_controller.py:973" *)
  wire \$465 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$467 ;
  (* src = "sdram_controller.py:399" *)
  wire \$469 ;
  (* src = "sdram_controller.py:727" *)
  wire \$47 ;
  (* src = "sdram_controller.py:400" *)
  wire \$471 ;
  (* src = "sdram_controller.py:399" *)
  wire \$473 ;
  (* src = "sdram_controller.py:403" *)
  wire \$475 ;
  (* src = "sdram_controller.py:406" *)
  wire \$477 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$479 ;
  (* src = "sdram_controller.py:1022" *)
  wire \$481 ;
  (* src = "sdram_controller.py:537" *)
  wire \$483 ;
  (* src = "sdram_controller.py:540" *)
  wire \$485 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$487 ;
  (* src = "sdram_controller.py:613" *)
  wire \$489 ;
  (* src = "sdram_controller.py:773" *)
  wire \$49 ;
  (* src = "sdram_controller.py:614" *)
  wire \$491 ;
  (* src = "sdram_controller.py:613" *)
  wire \$493 ;
  (* src = "sdram_controller.py:617" *)
  wire \$495 ;
  (* src = "sdram_controller.py:620" *)
  wire \$497 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$499 ;
  (* src = "sdram_controller.py:659" *)
  wire \$5 ;
  (* src = "sdram_controller.py:537" *)
  wire \$501 ;
  (* src = "sdram_controller.py:540" *)
  wire \$503 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$505 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$507 ;
  (* src = "sdram_controller.py:356" *)
  wire \$509 ;
  (* src = "sdram_controller.py:801" *)
  wire \$51 ;
  (* src = "sdram_controller.py:359" *)
  wire \$511 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$513 ;
  (* src = "sdram_controller.py:537" *)
  wire \$515 ;
  (* src = "sdram_controller.py:540" *)
  wire \$517 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$519 ;
  (* src = "sdram_controller.py:547" *)
  wire \$521 ;
  (* src = "sdram_controller.py:550" *)
  wire \$523 ;
  (* src = "sdram_controller.py:553" *)
  wire \$525 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$527 ;
  (* src = "sdram_controller.py:537" *)
  wire \$529 ;
  (* src = "sdram_controller.py:824" *)
  wire \$53 ;
  (* src = "sdram_controller.py:540" *)
  wire \$531 ;
  (* src = "sdram_controller.py:716" *)
  wire \$533 ;
  (* src = "sdram_controller.py:540" *)
  wire \$535 ;
  (* src = "sdram_controller.py:741" *)
  wire \$537 ;
  (* src = "sdram_controller.py:390" *)
  wire \$539 ;
  (* src = "sdram_controller.py:392" *)
  wire \$541 ;
  (* src = "sdram_controller.py:746" *)
  wire \$543 ;
  (* src = "sdram_controller.py:540" *)
  wire \$545 ;
  (* src = "sdram_controller.py:750" *)
  wire \$547 ;
  (* src = "sdram_controller.py:487" *)
  wire \$549 ;
  (* src = "sdram_controller.py:958" *)
  wire \$55 ;
  (* src = "sdram_controller.py:501" *)
  wire \$551 ;
  (* src = "sdram_controller.py:503" *)
  wire \$553 ;
  (* src = "sdram_controller.py:758" *)
  wire \$555 ;
  (* src = "sdram_controller.py:547" *)
  wire \$557 ;
  (* src = "sdram_controller.py:553" *)
  wire \$559 ;
  (* src = "sdram_controller.py:762" *)
  wire \$561 ;
  (* src = "sdram_controller.py:540" *)
  wire \$563 ;
  (* src = "sdram_controller.py:512" *)
  wire \$565 ;
  (* src = "sdram_controller.py:824" *)
  wire \$567 ;
  (* src = "sdram_controller.py:329" *)
  wire \$569 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$57 ;
  (* src = "sdram_controller.py:329" *)
  wire \$571 ;
  (* src = "sdram_controller.py:329" *)
  wire \$573 ;
  (* src = "sdram_controller.py:331" *)
  wire \$575 ;
  (* src = "sdram_controller.py:334" *)
  wire \$577 ;
  (* src = "sdram_controller.py:834" *)
  wire \$579 ;
  (* src = "sdram_controller.py:540" *)
  wire \$581 ;
  (* src = "sdram_controller.py:840" *)
  wire \$583 ;
  (* src = "sdram_controller.py:841" *)
  wire \$585 ;
  (* src = "sdram_controller.py:843" *)
  wire \$587 ;
  (* src = "sdram_controller.py:443" *)
  wire \$589 ;
  (* src = "sdram_controller.py:1103" *)
  wire \$59 ;
  (* src = "sdram_controller.py:444" *)
  wire \$591 ;
  (* src = "sdram_controller.py:443" *)
  wire \$593 ;
  (* src = "sdram_controller.py:450" *)
  wire \$595 ;
  (* src = "sdram_controller.py:853" *)
  wire \$597 ;
  (* src = "sdram_controller.py:540" *)
  wire \$599 ;
  (* src = "sdram_controller.py:872" *)
  wire \$601 ;
  (* src = "sdram_controller.py:918" *)
  wire \$603 ;
  (* src = "sdram_controller.py:613" *)
  wire \$605 ;
  (* src = "sdram_controller.py:614" *)
  wire \$607 ;
  (* src = "sdram_controller.py:613" *)
  wire \$609 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$61 ;
  (* src = "sdram_controller.py:620" *)
  wire \$611 ;
  (* src = "sdram_controller.py:920" *)
  wire \$613 ;
  (* src = "sdram_controller.py:359" *)
  wire \$615 ;
  (* src = "sdram_controller.py:929" *)
  wire \$617 ;
  (* src = "sdram_controller.py:540" *)
  wire \$619 ;
  (* src = "sdram_controller.py:958" *)
  wire \$621 ;
  (* src = "sdram_controller.py:329" *)
  wire \$623 ;
  (* src = "sdram_controller.py:329" *)
  wire \$625 ;
  (* src = "sdram_controller.py:329" *)
  wire \$627 ;
  (* src = "sdram_controller.py:331" *)
  wire \$629 ;
  (* src = "sdram_controller.py:1105" *)
  wire \$63 ;
  (* src = "sdram_controller.py:334" *)
  wire \$631 ;
  (* src = "sdram_controller.py:967" *)
  wire \$633 ;
  (* src = "sdram_controller.py:540" *)
  wire \$635 ;
  (* src = "sdram_controller.py:973" *)
  wire \$637 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$639 ;
  (* src = "sdram_controller.py:399" *)
  wire \$641 ;
  (* src = "sdram_controller.py:400" *)
  wire \$643 ;
  (* src = "sdram_controller.py:399" *)
  wire \$645 ;
  (* src = "sdram_controller.py:406" *)
  wire \$647 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$649 ;
  (* src = "sdram_controller.py:716" *)
  wire \$65 ;
  (* src = "sdram_controller.py:1022" *)
  wire \$651 ;
  (* src = "sdram_controller.py:540" *)
  wire \$653 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$655 ;
  (* src = "sdram_controller.py:613" *)
  wire \$657 ;
  (* src = "sdram_controller.py:614" *)
  wire \$659 ;
  (* src = "sdram_controller.py:613" *)
  wire \$661 ;
  (* src = "sdram_controller.py:620" *)
  wire \$663 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$665 ;
  (* src = "sdram_controller.py:540" *)
  wire \$667 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$669 ;
  (* src = "sdram_controller.py:741" *)
  wire \$67 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$671 ;
  (* src = "sdram_controller.py:359" *)
  wire \$673 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$675 ;
  (* src = "sdram_controller.py:540" *)
  wire \$677 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$679 ;
  (* src = "sdram_controller.py:547" *)
  wire \$681 ;
  (* src = "sdram_controller.py:553" *)
  wire \$683 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$685 ;
  (* src = "sdram_controller.py:540" *)
  wire \$687 ;
  (* src = "sdram_controller.py:716" *)
  wire \$689 ;
  (* src = "sdram_controller.py:746" *)
  wire \$69 ;
  (* src = "sdram_controller.py:540" *)
  wire \$691 ;
  (* src = "sdram_controller.py:741" *)
  wire \$693 ;
  (* src = "sdram_controller.py:378" *)
  wire \$695 ;
  (* src = "sdram_controller.py:746" *)
  wire \$697 ;
  (* src = "sdram_controller.py:540" *)
  wire \$699 ;
  (* src = "sdram_controller.py:659" *)
  wire \$7 ;
  (* src = "sdram_controller.py:750" *)
  wire \$701 ;
  (* src = "sdram_controller.py:487" *)
  wire \$703 ;
  (* src = "sdram_controller.py:493" *)
  wire \$705 ;
  (* src = "sdram_controller.py:758" *)
  wire \$707 ;
  (* src = "sdram_controller.py:547" *)
  wire \$709 ;
  (* src = "sdram_controller.py:750" *)
  wire \$71 ;
  (* src = "sdram_controller.py:553" *)
  wire \$711 ;
  (* src = "sdram_controller.py:762" *)
  wire \$713 ;
  (* src = "sdram_controller.py:540" *)
  wire \$715 ;
  (* src = "sdram_controller.py:512" *)
  wire \$717 ;
  (* src = "sdram_controller.py:824" *)
  wire \$719 ;
  (* src = "sdram_controller.py:329" *)
  wire \$721 ;
  (* src = "sdram_controller.py:329" *)
  wire \$723 ;
  (* src = "sdram_controller.py:329" *)
  wire \$725 ;
  (* src = "sdram_controller.py:331" *)
  wire \$727 ;
  (* src = "sdram_controller.py:334" *)
  wire \$729 ;
  (* src = "sdram_controller.py:758" *)
  wire \$73 ;
  (* src = "sdram_controller.py:834" *)
  wire \$731 ;
  (* src = "sdram_controller.py:540" *)
  wire \$733 ;
  (* src = "sdram_controller.py:840" *)
  wire \$735 ;
  (* src = "sdram_controller.py:841" *)
  wire \$737 ;
  (* src = "sdram_controller.py:843" *)
  wire \$739 ;
  (* src = "sdram_controller.py:443" *)
  wire \$741 ;
  (* src = "sdram_controller.py:444" *)
  wire \$743 ;
  (* src = "sdram_controller.py:443" *)
  wire \$745 ;
  (* src = "sdram_controller.py:450" *)
  wire \$747 ;
  (* src = "sdram_controller.py:853" *)
  wire \$749 ;
  (* src = "sdram_controller.py:762" *)
  wire \$75 ;
  (* src = "sdram_controller.py:540" *)
  wire \$751 ;
  (* src = "sdram_controller.py:920" *)
  wire \$753 ;
  (* src = "sdram_controller.py:359" *)
  wire \$755 ;
  (* src = "sdram_controller.py:929" *)
  wire \$757 ;
  (* src = "sdram_controller.py:540" *)
  wire \$759 ;
  (* src = "sdram_controller.py:958" *)
  wire \$761 ;
  (* src = "sdram_controller.py:329" *)
  wire \$763 ;
  (* src = "sdram_controller.py:329" *)
  wire \$765 ;
  (* src = "sdram_controller.py:329" *)
  wire \$767 ;
  (* src = "sdram_controller.py:331" *)
  wire \$769 ;
  (* src = "sdram_controller.py:824" *)
  wire \$77 ;
  (* src = "sdram_controller.py:334" *)
  wire \$771 ;
  (* src = "sdram_controller.py:967" *)
  wire \$773 ;
  (* src = "sdram_controller.py:540" *)
  wire \$775 ;
  (* src = "sdram_controller.py:973" *)
  wire \$777 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$779 ;
  (* src = "sdram_controller.py:399" *)
  wire \$781 ;
  (* src = "sdram_controller.py:400" *)
  wire \$783 ;
  (* src = "sdram_controller.py:399" *)
  wire \$785 ;
  (* src = "sdram_controller.py:406" *)
  wire \$787 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$789 ;
  (* src = "sdram_controller.py:834" *)
  wire \$79 ;
  (* src = "sdram_controller.py:1022" *)
  wire \$791 ;
  (* src = "sdram_controller.py:540" *)
  wire \$793 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$795 ;
  (* src = "sdram_controller.py:540" *)
  wire \$797 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$799 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$801 ;
  (* src = "sdram_controller.py:359" *)
  wire \$803 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$805 ;
  (* src = "sdram_controller.py:540" *)
  wire \$807 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$809 ;
  (* src = "sdram_controller.py:840" *)
  wire \$81 ;
  (* src = "sdram_controller.py:547" *)
  wire \$811 ;
  (* src = "sdram_controller.py:553" *)
  wire \$813 ;
  (* src = "sdram_controller.py:1101" *)
  wire \$815 ;
  (* src = "sdram_controller.py:540" *)
  wire \$817 ;
  (* src = "sdram_controller.py:716" *)
  wire \$819 ;
  (* src = "sdram_controller.py:741" *)
  wire \$821 ;
  (* src = "sdram_controller.py:773" *)
  wire \$823 ;
  (* src = "sdram_controller.py:716" *)
  wire \$825 ;
  (* src = "sdram_controller.py:726" *)
  wire \$827 ;
  (* src = "sdram_controller.py:727" *)
  wire \$829 ;
  (* src = "sdram_controller.py:841" *)
  wire \$83 ;
  (* src = "sdram_controller.py:728" *)
  wire [15:0] \$831 ;
  (* src = "sdram_controller.py:728" *)
  wire [15:0] \$832 ;
  (* src = "sdram_controller.py:716" *)
  wire \$834 ;
  (* src = "sdram_controller.py:726" *)
  wire \$836 ;
  (* src = "sdram_controller.py:727" *)
  wire \$838 ;
  (* src = "sdram_controller.py:741" *)
  wire \$840 ;
  (* src = "sdram_controller.py:746" *)
  wire \$842 ;
  (* src = "sdram_controller.py:750" *)
  wire \$844 ;
  (* src = "sdram_controller.py:758" *)
  wire \$846 ;
  (* src = "sdram_controller.py:762" *)
  wire \$848 ;
  (* src = "sdram_controller.py:843" *)
  wire \$85 ;
  (* src = "sdram_controller.py:767" *)
  wire \$850 ;
  (* src = "sdram_controller.py:768" *)
  wire \$852 ;
  (* src = "sdram_controller.py:770" *)
  wire \$854 ;
  (* src = "sdram_controller.py:773" *)
  wire \$856 ;
  (* src = "sdram_controller.py:818" *)
  wire \$858 ;
  (* src = "sdram_controller.py:824" *)
  wire \$860 ;
  (* src = "sdram_controller.py:834" *)
  wire \$862 ;
  (* src = "sdram_controller.py:840" *)
  wire \$864 ;
  (* src = "sdram_controller.py:841" *)
  wire \$866 ;
  (* src = "sdram_controller.py:843" *)
  wire \$868 ;
  (* src = "sdram_controller.py:853" *)
  wire \$87 ;
  (* src = "sdram_controller.py:853" *)
  wire \$870 ;
  (* src = "sdram_controller.py:858" *)
  wire \$872 ;
  (* src = "sdram_controller.py:866" *)
  wire \$874 ;
  (* src = "sdram_controller.py:872" *)
  wire \$876 ;
  (* src = "sdram_controller.py:913" *)
  wire \$878 ;
  (* src = "sdram_controller.py:920" *)
  wire \$880 ;
  (* src = "sdram_controller.py:929" *)
  wire \$882 ;
  (* src = "sdram_controller.py:935" *)
  wire \$884 ;
  (* src = "sdram_controller.py:939" *)
  wire \$886 ;
  (* src = "sdram_controller.py:954" *)
  wire \$888 ;
  (* src = "sdram_controller.py:872" *)
  wire \$89 ;
  (* src = "sdram_controller.py:958" *)
  wire \$890 ;
  (* src = "sdram_controller.py:967" *)
  wire \$892 ;
  (* src = "sdram_controller.py:973" *)
  wire \$894 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$896 ;
  (* src = "sdram_controller.py:1015" *)
  wire \$898 ;
  (* src = "sdram_controller.py:726" *)
  wire \$9 ;
  (* src = "sdram_controller.py:1054" *)
  wire \$900 ;
  (* src = "sdram_controller.py:1065" *)
  wire \$902 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$904 ;
  (* src = "sdram_controller.py:1080" *)
  wire \$906 ;
  (* src = "sdram_controller.py:1084" *)
  wire \$908 ;
  (* src = "sdram_controller.py:918" *)
  wire \$91 ;
  (* src = "sdram_controller.py:716" *)
  wire \$910 ;
  (* src = "sdram_controller.py:741" *)
  wire \$912 ;
  (* src = "sdram_controller.py:378" *)
  wire \$914 ;
  (* src = "sdram_controller.py:750" *)
  wire \$916 ;
  (* src = "sdram_controller.py:487" *)
  wire \$918 ;
  (* src = "sdram_controller.py:493" *)
  wire \$920 ;
  (* src = "sdram_controller.py:758" *)
  wire \$922 ;
  (* src = "sdram_controller.py:547" *)
  wire \$924 ;
  (* src = "sdram_controller.py:553" *)
  wire \$926 ;
  (* src = "sdram_controller.py:512" *)
  wire \$928 ;
  (* src = "sdram_controller.py:920" *)
  wire \$93 ;
  (* src = "sdram_controller.py:824" *)
  wire \$930 ;
  (* src = "sdram_controller.py:329" *)
  wire \$932 ;
  (* src = "sdram_controller.py:329" *)
  wire \$934 ;
  (* src = "sdram_controller.py:329" *)
  wire \$936 ;
  (* src = "sdram_controller.py:331" *)
  wire \$938 ;
  (* src = "sdram_controller.py:334" *)
  wire \$940 ;
  (* src = "sdram_controller.py:840" *)
  wire \$942 ;
  (* src = "sdram_controller.py:841" *)
  wire \$944 ;
  (* src = "sdram_controller.py:843" *)
  wire \$946 ;
  (* src = "sdram_controller.py:443" *)
  wire \$948 ;
  (* src = "sdram_controller.py:929" *)
  wire \$95 ;
  (* src = "sdram_controller.py:444" *)
  wire \$950 ;
  (* src = "sdram_controller.py:443" *)
  wire \$952 ;
  (* src = "sdram_controller.py:450" *)
  wire \$954 ;
  (* src = "sdram_controller.py:920" *)
  wire \$956 ;
  (* src = "sdram_controller.py:359" *)
  wire \$958 ;
  (* src = "sdram_controller.py:958" *)
  wire \$960 ;
  (* src = "sdram_controller.py:329" *)
  wire \$962 ;
  (* src = "sdram_controller.py:329" *)
  wire \$964 ;
  (* src = "sdram_controller.py:329" *)
  wire \$966 ;
  (* src = "sdram_controller.py:331" *)
  wire \$968 ;
  (* src = "sdram_controller.py:958" *)
  wire \$97 ;
  (* src = "sdram_controller.py:334" *)
  wire \$970 ;
  (* src = "sdram_controller.py:973" *)
  wire \$972 ;
  (* src = "sdram_controller.py:1002" *)
  wire \$974 ;
  (* src = "sdram_controller.py:399" *)
  wire \$976 ;
  (* src = "sdram_controller.py:400" *)
  wire \$978 ;
  (* src = "sdram_controller.py:399" *)
  wire \$980 ;
  (* src = "sdram_controller.py:406" *)
  wire \$982 ;
  (* src = "sdram_controller.py:1071" *)
  wire \$984 ;
  (* src = "sdram_controller.py:1074" *)
  wire \$986 ;
  (* src = "sdram_controller.py:359" *)
  wire \$988 ;
  (* src = "sdram_controller.py:967" *)
  wire \$99 ;
  (* src = "sdram_controller.py:1096" *)
  wire \$990 ;
  (* src = "sdram_controller.py:547" *)
  wire \$992 ;
  (* src = "sdram_controller.py:553" *)
  wire \$994 ;
  (* src = "sdram_controller.py:716" *)
  wire \$996 ;
  (* src = "sdram_controller.py:741" *)
  wire \$998 ;
  (* src = "sdram_controller.py:239" *)
  reg allBanksIdle;
  (* src = "sdram_controller.py:1179" *)
  reg bankController0_bankActivated;
  (* src = "sdram_controller.py:1178" *)
  wire bankController0_bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  wire bankController0_bankCanPreCharge;
  (* src = "sdram_controller.py:1171" *)
  wire [9:0] bankController0_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1176" *)
  wire bankController0_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] bankController0_bankState = 3'h0;
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] \bankController0_bankState$next ;
  (* src = "sdram_controller.py:1180" *)
  reg bankController0_otherBankActivated;
  (* src = "sdram_controller.py:1179" *)
  reg bankController1_bankActivated;
  (* src = "sdram_controller.py:1178" *)
  wire bankController1_bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  wire bankController1_bankCanPreCharge;
  (* src = "sdram_controller.py:1171" *)
  wire [9:0] bankController1_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1176" *)
  wire bankController1_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] bankController1_bankState = 3'h0;
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] \bankController1_bankState$next ;
  (* src = "sdram_controller.py:1180" *)
  reg bankController1_otherBankActivated;
  (* src = "sdram_controller.py:1179" *)
  reg bankController2_bankActivated;
  (* src = "sdram_controller.py:1178" *)
  wire bankController2_bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  wire bankController2_bankCanPreCharge;
  (* src = "sdram_controller.py:1171" *)
  wire [9:0] bankController2_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1176" *)
  wire bankController2_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] bankController2_bankState = 3'h0;
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] \bankController2_bankState$next ;
  (* src = "sdram_controller.py:1180" *)
  reg bankController2_otherBankActivated;
  (* src = "sdram_controller.py:1179" *)
  reg bankController3_bankActivated;
  (* src = "sdram_controller.py:1178" *)
  wire bankController3_bankCanActivate;
  (* src = "sdram_controller.py:1177" *)
  wire bankController3_bankCanPreCharge;
  (* src = "sdram_controller.py:1171" *)
  wire [9:0] bankController3_bankREFIcyclesCounter;
  (* src = "sdram_controller.py:1176" *)
  wire bankController3_bankShouldRefresh;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] bankController3_bankState = 3'h0;
  (* src = "sdram_controller.py:1175" *)
  reg [2:0] \bankController3_bankState$next ;
  (* src = "sdram_controller.py:1180" *)
  reg bankController3_otherBankActivated;
  (* src = "sdram_controller.py:238" *)
  reg banksShouldRefresh;
  (* src = "sdram_controller.py:261" *)
  reg burstWritesMode = 1'h0;
  (* src = "sdram_controller.py:261" *)
  reg \burstWritesMode$next ;
  (* src = "sdram_controller.py:1290" *)
  wire clkSDRAM_clk;
  (* src = "sdram_controller.py:1290" *)
  wire clkSDRAM_rst;
  (* src = "sdram_controller.py:254" *)
  reg cmdCompleted;
  (* src = "sdram_controller.py:255" *)
  reg [3:0] cmdIndex = 4'h0;
  (* src = "sdram_controller.py:255" *)
  reg [3:0] \cmdIndex$next ;
  (* src = "sdram_controller.py:253" *)
  reg [1:0] cmdRemainingCyclesCounter;
  (* src = "sdram_controller.py:249" *)
  reg [20:0] ctrlAddress = 21'h000000;
  (* src = "sdram_controller.py:249" *)
  reg [20:0] \ctrlAddress$next ;
  (* src = "sdram_controller.py:222" *)
  input ctrlRd;
  wire ctrlRd;
  (* src = "sdram_controller.py:221" *)
  input [20:0] ctrlRdAddress;
  wire [20:0] ctrlRdAddress;
  (* src = "sdram_controller.py:223" *)
  output [23:0] ctrlRdDataOut;
  reg [23:0] ctrlRdDataOut;
  (* src = "sdram_controller.py:225" *)
  reg ctrlRdInProgress = 1'h0;
  (* src = "sdram_controller.py:225" *)
  reg \ctrlRdInProgress$next ;
  (* src = "sdram_controller.py:224" *)
  output ctrlRdIncAddress;
  reg ctrlRdIncAddress = 1'h0;
  (* src = "sdram_controller.py:224" *)
  reg \ctrlRdIncAddress$next ;
  (* src = "sdram_controller.py:213" *)
  output ctrlReady;
  reg ctrlReady = 1'h0;
  (* src = "sdram_controller.py:213" *)
  reg \ctrlReady$next ;
  (* src = "sdram_controller.py:216" *)
  input ctrlWr;
  wire ctrlWr;
  (* src = "sdram_controller.py:215" *)
  input [20:0] ctrlWrAddress;
  wire [20:0] ctrlWrAddress;
  (* src = "sdram_controller.py:217" *)
  input [23:0] ctrlWrDataIn;
  wire [23:0] ctrlWrDataIn;
  (* src = "sdram_controller.py:219" *)
  reg ctrlWrInProgress = 1'h0;
  (* src = "sdram_controller.py:219" *)
  reg \ctrlWrInProgress$next ;
  (* src = "sdram_controller.py:218" *)
  output ctrlWrIncAddress;
  reg ctrlWrIncAddress = 1'h0;
  (* src = "sdram_controller.py:218" *)
  reg \ctrlWrIncAddress$next ;
  (* enum_base_type = "Command" *)
  (* enum_value_00000 = "NoCommand" *)
  (* enum_value_00001 = "BankActivate" *)
  (* enum_value_00010 = "BankPreCharge" *)
  (* enum_value_00011 = "PreChargeAll" *)
  (* enum_value_00100 = "Write" *)
  (* enum_value_00101 = "WriteAndAutoPreCharge" *)
  (* enum_value_00110 = "Read" *)
  (* enum_value_00111 = "ReadAndAutoPreCharge" *)
  (* enum_value_01000 = "ModeRegisterSet" *)
  (* enum_value_01001 = "NoOperation" *)
  (* enum_value_01010 = "BurstStop" *)
  (* enum_value_01011 = "DeviceDeSelect" *)
  (* enum_value_01100 = "AutoRefresh" *)
  (* enum_value_01101 = "SelfRefreshEntry" *)
  (* enum_value_01110 = "SelfRefreshExit" *)
  (* enum_value_01111 = "ClockSuspendModeExit" *)
  (* enum_value_10000 = "PowerDownModeExit" *)
  (* enum_value_10001 = "DataWrite_OutputEnable" *)
  (* enum_value_10010 = "DataMask_OutputDisable" *)
  (* src = "sdram_controller.py:252" *)
  reg [4:0] currentCommand = 5'h00;
  (* src = "sdram_controller.py:252" *)
  reg [4:0] \currentCommand$next ;
  (* enum_base_type = "SDRAMControllerStates" *)
  (* enum_value_000 = "InitOp" *)
  (* enum_value_001 = "ConfigurationOp" *)
  (* enum_value_010 = "Idle" *)
  (* enum_value_011 = "RefreshOp" *)
  (* enum_value_100 = "WriteBurstOp" *)
  (* enum_value_101 = "WriteOp" *)
  (* enum_value_110 = "ReadOp" *)
  (* enum_value_111 = "Error" *)
  (* src = "sdram_controller.py:230" *)
  reg [2:0] currentControllerState;
  (* src = "sdram_controller.py:259" *)
  reg [4:0] delayCounter = 5'h00;
  (* src = "sdram_controller.py:259" *)
  reg [4:0] \delayCounter$next ;
  (* src = "sdram_controller.py:228" *)
  reg errorState = 1'h0;
  (* src = "sdram_controller.py:228" *)
  reg \errorState$next ;
  (* enum_base_type = "Command" *)
  (* enum_value_00000 = "NoCommand" *)
  (* enum_value_00001 = "BankActivate" *)
  (* enum_value_00010 = "BankPreCharge" *)
  (* enum_value_00011 = "PreChargeAll" *)
  (* enum_value_00100 = "Write" *)
  (* enum_value_00101 = "WriteAndAutoPreCharge" *)
  (* enum_value_00110 = "Read" *)
  (* enum_value_00111 = "ReadAndAutoPreCharge" *)
  (* enum_value_01000 = "ModeRegisterSet" *)
  (* enum_value_01001 = "NoOperation" *)
  (* enum_value_01010 = "BurstStop" *)
  (* enum_value_01011 = "DeviceDeSelect" *)
  (* enum_value_01100 = "AutoRefresh" *)
  (* enum_value_01101 = "SelfRefreshEntry" *)
  (* enum_value_01110 = "SelfRefreshExit" *)
  (* enum_value_01111 = "ClockSuspendModeExit" *)
  (* enum_value_10000 = "PowerDownModeExit" *)
  (* enum_value_10001 = "DataWrite_OutputEnable" *)
  (* enum_value_10010 = "DataMask_OutputDisable" *)
  (* src = "sdram_controller.py:251" *)
  reg [4:0] nextCommand;
  (* src = "sdram_controller.py:262" *)
  reg [7:0] pageColumnIndex = 8'h00;
  (* src = "sdram_controller.py:262" *)
  reg [7:0] \pageColumnIndex$next ;
  (* src = "sdram_controller.py:258" *)
  reg [14:0] powerUpCounter = 15'h0000;
  (* src = "sdram_controller.py:258" *)
  reg [14:0] \powerUpCounter$next ;
  (* enum_base_type = "SDRAMControllerStates" *)
  (* enum_value_000 = "InitOp" *)
  (* enum_value_001 = "ConfigurationOp" *)
  (* enum_value_010 = "Idle" *)
  (* enum_value_011 = "RefreshOp" *)
  (* enum_value_100 = "WriteBurstOp" *)
  (* enum_value_101 = "WriteOp" *)
  (* enum_value_110 = "ReadOp" *)
  (* enum_value_111 = "Error" *)
  (* src = "sdram_controller.py:231" *)
  reg [2:0] previousControllerState = 3'h0;
  (* src = "sdram_controller.py:231" *)
  reg [2:0] \previousControllerState$next ;
  (* src = "sdram_controller.py:256" *)
  reg refreshCmdIndex = 1'h0;
  (* src = "sdram_controller.py:256" *)
  reg \refreshCmdIndex$next ;
  (* src = "sdram_controller.py:257" *)
  reg refreshRequired = 1'h0;
  (* src = "sdram_controller.py:257" *)
  reg \refreshRequired$next ;
  (* src = "sdram_controller.py:706" *)
  reg repeatRefresh = 1'h0;
  (* src = "sdram_controller.py:706" *)
  reg \repeatRefresh$next ;
  (* src = "sdram_controller.py:205" *)
  output [10:0] sdramAddress;
  reg [10:0] sdramAddress = 11'h000;
  (* src = "sdram_controller.py:205" *)
  reg [10:0] \sdramAddress$next ;
  (* src = "sdram_controller.py:206" *)
  output [1:0] sdramBank;
  reg [1:0] sdramBank = 2'h0;
  (* src = "sdram_controller.py:206" *)
  reg [1:0] \sdramBank$next ;
  (* src = "sdram_controller.py:202" *)
  output sdramCASn;
  reg sdramCASn = 1'h0;
  (* src = "sdram_controller.py:202" *)
  reg \sdramCASn$next ;
  (* src = "sdram_controller.py:204" *)
  output sdramCSn;
  reg sdramCSn = 1'h0;
  (* src = "sdram_controller.py:204" *)
  reg \sdramCSn$next ;
  (* src = "sdram_controller.py:199" *)
  output sdramClk;
  wire sdramClk;
  (* src = "sdram_controller.py:200" *)
  output sdramClkEn;
  reg sdramClkEn = 1'h0;
  (* src = "sdram_controller.py:200" *)
  reg \sdramClkEn$next ;
  (* src = "sdram_controller.py:708" *)
  reg [2:0] sdramCtrlr_state = 3'h0;
  (* src = "sdram_controller.py:708" *)
  reg [2:0] \sdramCtrlr_state$next ;
  (* src = "sdram_controller.py:210" *)
  output [3:0] sdramDataMasks;
  reg [3:0] sdramDataMasks = 4'hf;
  (* src = "sdram_controller.py:210" *)
  reg [3:0] \sdramDataMasks$next ;
  (* src = "sdram_controller.py:208" *)
  output [31:0] sdramDqIn;
  reg [31:0] sdramDqIn = 32'd0;
  (* src = "sdram_controller.py:208" *)
  reg [31:0] \sdramDqIn$next ;
  (* src = "sdram_controller.py:207" *)
  input [31:0] sdramDqOut;
  wire [31:0] sdramDqOut;
  (* src = "sdram_controller.py:209" *)
  output sdramDqWRn;
  reg sdramDqWRn = 1'h0;
  (* src = "sdram_controller.py:209" *)
  reg \sdramDqWRn$next ;
  (* src = "sdram_controller.py:201" *)
  output sdramRASn;
  reg sdramRASn = 1'h0;
  (* src = "sdram_controller.py:201" *)
  reg \sdramRASn$next ;
  (* src = "sdram_controller.py:203" *)
  output sdramWEn;
  reg sdramWEn = 1'h0;
  (* src = "sdram_controller.py:203" *)
  reg \sdramWEn$next ;
  (* src = "sdram_controller.py:233" *)
  wire [1:0] targetBankAddress;
  (* src = "sdram_controller.py:240" *)
  reg targetBankCanActivate = 1'h0;
  (* src = "sdram_controller.py:240" *)
  reg \targetBankCanActivate$next ;
  (* src = "sdram_controller.py:241" *)
  reg targetBankCanPreCharge = 1'h0;
  (* src = "sdram_controller.py:241" *)
  reg \targetBankCanPreCharge$next ;
  (* src = "sdram_controller.py:242" *)
  reg [9:0] targetBankRefreshCounter = 10'h000;
  (* src = "sdram_controller.py:242" *)
  reg [9:0] \targetBankRefreshCounter$next ;
  (* enum_base_type = "BankControllerStates" *)
  (* enum_value_000 = "NotReady" *)
  (* enum_value_001 = "Idle" *)
  (* enum_value_010 = "Active" *)
  (* enum_value_011 = "ActiveBurst" *)
  (* enum_value_100 = "PreCharge" *)
  (* enum_value_101 = "Refreshing" *)
  (* src = "sdram_controller.py:243" *)
  reg [2:0] targetBankState;
  (* src = "sdram_controller.py:235" *)
  wire [7:0] targetColumnAddress;
  (* src = "sdram_controller.py:236" *)
  wire [3:0] targetMask;
  (* src = "sdram_controller.py:234" *)
  wire [10:0] targetRowAddress;
  assign \$9  = cmdIndex == (* src = "sdram_controller.py:726" *) 1'h1;
  assign \$99  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$1002  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1004  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$1008  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1010  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1016  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1018  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$101  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1020  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1022  = \$1018  | (* src = "sdram_controller.py:329" *) \$1020 ;
  assign \$1024  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1028  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1030  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$1032  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$1034  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$1036  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$1038  = \$1034  & (* src = "sdram_controller.py:443" *) \$1036 ;
  assign \$103  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$1042  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$1046  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1048  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1050  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1052  = \$1048  | (* src = "sdram_controller.py:329" *) \$1050 ;
  assign \$1054  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1058  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$105  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$1060  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$1062  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$1064  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$1066  = \$1062  & (* src = "sdram_controller.py:399" *) \$1064 ;
  assign \$1070  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1072  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1076  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1078  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$107  = pageColumnIndex == (* src = "sdram_controller.py:1022" *) targetColumnAddress;
  assign \$1082  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$1084  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1088  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1090  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$1094  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1096  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$109  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$1102  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1104  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1106  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1108  = \$1104  | (* src = "sdram_controller.py:329" *) \$1106 ;
  assign \$1110  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1114  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1116  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$1118  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$111  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$1120  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$1122  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$1124  = \$1120  & (* src = "sdram_controller.py:443" *) \$1122 ;
  assign \$1128  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$1132  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1134  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1136  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1138  = \$1134  | (* src = "sdram_controller.py:329" *) \$1136 ;
  assign \$113  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1140  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1144  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1146  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$1148  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$1150  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$1152  = \$1148  & (* src = "sdram_controller.py:399" *) \$1150 ;
  assign \$1156  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1158  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$115  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1162  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1164  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1168  = cmdIndex == (* src = "sdram_controller.py:726" *) 1'h1;
  assign \$1170  = powerUpCounter > (* src = "sdram_controller.py:727" *) 1'h0;
  assign \$1172  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1176  = $signed(delayCounter) > (* src = "sdram_controller.py:390" *) $signed(5'h00);
  assign \$1178  = ! (* src = "sdram_controller.py:392" *) $signed(delayCounter);
  assign \$117  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$1181  = $signed(delayCounter) - (* src = "sdram_controller.py:391" *) $signed(5'h01);
  assign \$1183  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1185  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$1189  = $signed(delayCounter) > (* src = "sdram_controller.py:501" *) $signed(5'h00);
  assign \$1191  = ! (* src = "sdram_controller.py:503" *) $signed(delayCounter);
  assign \$1194  = $signed(delayCounter) - (* src = "sdram_controller.py:502" *) $signed(5'h01);
  assign \$1196  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$1198  = cmdIndex == (* src = "sdram_controller.py:767" *) 3'h5;
  assign \$11  = powerUpCounter > (* src = "sdram_controller.py:727" *) 1'h0;
  assign \$119  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1200  = $signed(delayCounter) > (* src = "sdram_controller.py:768" *) $signed(5'h00);
  assign \$1202  = ! (* src = "sdram_controller.py:770" *) $signed(delayCounter);
  assign \$1205  = $signed(delayCounter) - (* src = "sdram_controller.py:769" *) $signed(5'h01);
  assign \$1207  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$1209  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1211  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$1213  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$1216  = $signed(delayCounter) - (* src = "sdram_controller.py:842" *) $signed(5'h01);
  assign \$1218  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$1220  = cmdIndex == (* src = "sdram_controller.py:935" *) 4'ha;
  assign \$1222  = $signed(delayCounter) > (* src = "sdram_controller.py:937" *) $signed(5'h00);
  assign \$1225  = $signed(delayCounter) - (* src = "sdram_controller.py:938" *) $signed(5'h01);
  assign \$1227  = ! (* src = "sdram_controller.py:939" *) $signed(delayCounter);
  assign \$1229  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$1231  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1233  = $signed(delayCounter) > (* src = "sdram_controller.py:1000" *) $signed(5'h00);
  assign \$1236  = $signed(delayCounter) - (* src = "sdram_controller.py:1001" *) $signed(5'h01);
  assign \$1238  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$123  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$1240  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$1242  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$1244  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$1246  = $signed(delayCounter) > (* src = "sdram_controller.py:1067" *) $signed(5'h00);
  assign \$1249  = $signed(delayCounter) - (* src = "sdram_controller.py:1068" *) $signed(5'h01);
  assign \$1251  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1253  = $signed(delayCounter) > (* src = "sdram_controller.py:1072" *) $signed(5'h00);
  assign \$1256  = $signed(delayCounter) - (* src = "sdram_controller.py:1073" *) $signed(5'h01);
  assign \$1258  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$125  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1260  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$1262  = $signed(delayCounter) > (* src = "sdram_controller.py:1082" *) $signed(5'h00);
  assign \$1265  = $signed(delayCounter) - (* src = "sdram_controller.py:1083" *) $signed(5'h01);
  assign \$1267  = ! (* src = "sdram_controller.py:1084" *) $signed(delayCounter);
  assign \$1269  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1273  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$1275  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$1277  = \$1275  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$127  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$1280  = $signed(delayCounter) - (* src = "sdram_controller.py:1104" *) $signed(5'h01);
  assign \$1282  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1286  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1288  = ! (* src = "sdram_controller.py:752" *) cmdRemainingCyclesCounter;
  assign \$1290  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1292  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1294  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1296  = \$1292  | (* src = "sdram_controller.py:329" *) \$1294 ;
  assign \$1298  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$129  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1302  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1304  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$1306  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$1308  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$1310  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$1312  = \$1308  & (* src = "sdram_controller.py:443" *) \$1310 ;
  assign \$1316  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$131  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1320  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1322  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1324  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1326  = \$1322  | (* src = "sdram_controller.py:329" *) \$1324 ;
  assign \$1328  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1332  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1334  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$1336  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$1338  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$133  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$1340  = \$1336  & (* src = "sdram_controller.py:399" *) \$1338 ;
  assign \$1344  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1346  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1350  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1354  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1356  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$135  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1360  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$1362  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1364  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1366  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1368  = \$1364  | (* src = "sdram_controller.py:329" *) \$1366 ;
  assign \$1370  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1374  = ! (* src = "sdram_controller.py:338" *) targetBankAddress;
  assign \$1376  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$137  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$1380  = ! (* src = "sdram_controller.py:363" *) targetBankAddress;
  assign \$1382  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1384  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1386  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1388  = \$1384  | (* src = "sdram_controller.py:329" *) \$1386 ;
  assign \$1390  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1394  = ! (* src = "sdram_controller.py:338" *) targetBankAddress;
  assign \$1396  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1398  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$13  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$139  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1402  = ! (* src = "sdram_controller.py:363" *) targetBankAddress;
  assign \$1404  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1406  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1412  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$1414  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$1416  = \$1414  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$1418  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$141  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$1422  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1424  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1428  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$1430  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1432  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1434  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1436  = \$1432  | (* src = "sdram_controller.py:329" *) \$1434 ;
  assign \$1438  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$143  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$1442  = targetBankAddress == (* src = "sdram_controller.py:338" *) 1'h1;
  assign \$1444  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$1448  = targetBankAddress == (* src = "sdram_controller.py:363" *) 1'h1;
  assign \$1450  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1452  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1454  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1456  = \$1452  | (* src = "sdram_controller.py:329" *) \$1454 ;
  assign \$1458  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$145  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$1462  = targetBankAddress == (* src = "sdram_controller.py:338" *) 1'h1;
  assign \$1464  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1466  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1470  = targetBankAddress == (* src = "sdram_controller.py:363" *) 1'h1;
  assign \$1472  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1474  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$147  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$1480  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$1482  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$1484  = \$1482  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$1486  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1490  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1492  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1496  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$1498  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$149  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$1500  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1502  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1504  = \$1500  | (* src = "sdram_controller.py:329" *) \$1502 ;
  assign \$1506  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1510  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h2;
  assign \$1512  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$1516  = targetBankAddress == (* src = "sdram_controller.py:363" *) 2'h2;
  assign \$1518  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$151  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$1520  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1522  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1524  = \$1520  | (* src = "sdram_controller.py:329" *) \$1522 ;
  assign \$1526  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1530  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h2;
  assign \$1532  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1534  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1538  = targetBankAddress == (* src = "sdram_controller.py:363" *) 2'h2;
  assign \$153  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$1540  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1542  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1548  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$1550  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$1552  = \$1550  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$1554  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1558  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$155  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1560  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1564  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$1566  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1568  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1570  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1572  = \$1568  | (* src = "sdram_controller.py:329" *) \$1570 ;
  assign \$1574  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1578  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h3;
  assign \$157  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$1580  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$1584  = targetBankAddress == (* src = "sdram_controller.py:363" *) 2'h3;
  assign \$1586  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1588  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1590  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1592  = \$1588  | (* src = "sdram_controller.py:329" *) \$1590 ;
  assign \$1594  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1598  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h3;
  assign \$15  = ctrlWr & (* src = "sdram_controller.py:801" *) burstWritesMode;
  assign \$159  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1600  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1602  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1606  = targetBankAddress == (* src = "sdram_controller.py:363" *) 2'h3;
  assign \$1608  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1610  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1616  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$1618  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$161  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$1620  = \$1618  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$1622  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1624  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$1626  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$1628  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$1630  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1632  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1634  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1636  = \$1632  | (* src = "sdram_controller.py:329" *) \$1634 ;
  assign \$1638  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$163  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$1642  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1644  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$1646  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$1648  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$1650  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$1652  = \$1648  & (* src = "sdram_controller.py:443" *) \$1650 ;
  assign \$1654  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$1656  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$1658  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$165  = pageColumnIndex == (* src = "sdram_controller.py:1022" *) targetColumnAddress;
  assign \$1660  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$1662  = \$1658  & (* src = "sdram_controller.py:613" *) \$1660 ;
  assign \$1664  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1666  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1668  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1670  = \$1666  | (* src = "sdram_controller.py:329" *) \$1668 ;
  assign \$1672  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1676  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1678  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$167  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$1680  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$1682  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$1684  = \$1680  & (* src = "sdram_controller.py:399" *) \$1682 ;
  assign \$1686  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$1688  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$1690  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$1692  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$1694  = \$1690  & (* src = "sdram_controller.py:613" *) \$1692 ;
  assign \$1696  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1698  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$169  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$1700  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1702  = ! (* src = "sdram_controller.py:752" *) cmdRemainingCyclesCounter;
  assign \$1704  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1706  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1708  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1710  = \$1706  | (* src = "sdram_controller.py:329" *) \$1708 ;
  assign \$1712  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1716  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$1718  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$171  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$1720  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$1722  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$1724  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$1726  = \$1722  & (* src = "sdram_controller.py:443" *) \$1724 ;
  assign \$1730  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1732  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1734  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1736  = \$1732  | (* src = "sdram_controller.py:329" *) \$1734 ;
  assign \$1738  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$173  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$1742  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$1744  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$1746  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$1748  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$1750  = \$1746  & (* src = "sdram_controller.py:399" *) \$1748 ;
  assign \$1754  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1756  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$1758  = ctrlWr & (* src = "sdram_controller.py:801" *) burstWritesMode;
  assign \$175  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$1760  = cmdIndex == (* src = "sdram_controller.py:935" *) 4'ha;
  assign \$1762  = ! (* src = "sdram_controller.py:939" *) $signed(delayCounter);
  assign \$1764  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$1766  = ! (* src = "sdram_controller.py:1084" *) $signed(delayCounter);
  assign \$1768  = ctrlWr & (* src = "sdram_controller.py:801" *) burstWritesMode;
  assign \$1770  = ! (* src = "sdram_controller.py:818" *) cmdIndex;
  assign \$1772  = 9'h100 - (* src = "sdram_controller.py:822" *) targetColumnAddress;
  assign \$1776  = \$1774  + (* src = "sdram_controller.py:822" *) 4'hf;
  assign \$1778  = \$1776  + (* src = "sdram_controller.py:822" *) 3'h5;
  assign \$177  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$1780  = targetBankRefreshCounter < (* src = "sdram_controller.py:822" *) \$1778 ;
  assign \$1782  = ! (* src = "sdram_controller.py:954" *) cmdIndex;
  assign \$1784  = 9'h100 - (* src = "sdram_controller.py:956" *) targetColumnAddress;
  assign \$1788  = \$1786  + (* src = "sdram_controller.py:956" *) 4'hd;
  assign \$1790  = \$1788  + (* src = "sdram_controller.py:956" *) 3'h5;
  assign \$1792  = targetBankRefreshCounter < (* src = "sdram_controller.py:956" *) \$1790 ;
  assign \$1796  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$1798  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$17  = ~ (* src = "sdram_controller.py:799" *) ctrlReady;
  assign \$1800  = \$1798  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$1802  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1804  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1806  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1808  = \$1804  | (* src = "sdram_controller.py:329" *) \$1806 ;
  assign \$1810  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1814  = ! (* src = "sdram_controller.py:338" *) targetBankAddress;
  assign \$1816  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1818  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$181  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$1820  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1822  = \$1818  | (* src = "sdram_controller.py:329" *) \$1820 ;
  assign \$1824  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1828  = ! (* src = "sdram_controller.py:338" *) targetBankAddress;
  assign \$1830  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1832  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1834  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1836  = \$1832  | (* src = "sdram_controller.py:329" *) \$1834 ;
  assign \$1838  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$183  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$1842  = ! (* src = "sdram_controller.py:338" *) targetBankAddress;
  assign \$1844  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1846  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1848  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1850  = \$1846  | (* src = "sdram_controller.py:329" *) \$1848 ;
  assign \$1852  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1856  = ! (* src = "sdram_controller.py:338" *) targetBankAddress;
  assign \$1858  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$185  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$1860  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1862  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1864  = \$1860  | (* src = "sdram_controller.py:329" *) \$1862 ;
  assign \$1866  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1870  = targetBankAddress == (* src = "sdram_controller.py:338" *) 1'h1;
  assign \$1872  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1874  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1876  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1878  = \$1874  | (* src = "sdram_controller.py:329" *) \$1876 ;
  assign \$187  = ~ (* src = "sdram_controller.py:375" *) sdramClkEn;
  assign \$1880  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1884  = targetBankAddress == (* src = "sdram_controller.py:338" *) 1'h1;
  assign \$1886  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1888  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1890  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1892  = \$1888  | (* src = "sdram_controller.py:329" *) \$1890 ;
  assign \$1894  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1898  = targetBankAddress == (* src = "sdram_controller.py:338" *) 1'h1;
  assign \$189  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$1900  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1902  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1904  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1906  = \$1902  | (* src = "sdram_controller.py:329" *) \$1904 ;
  assign \$1908  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1912  = targetBankAddress == (* src = "sdram_controller.py:338" *) 1'h1;
  assign \$1914  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1916  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1918  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$191  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$1920  = \$1916  | (* src = "sdram_controller.py:329" *) \$1918 ;
  assign \$1922  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1926  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h2;
  assign \$1928  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1930  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1932  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1934  = \$1930  | (* src = "sdram_controller.py:329" *) \$1932 ;
  assign \$1936  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$193  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$1940  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h2;
  assign \$1942  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1944  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1946  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1948  = \$1944  | (* src = "sdram_controller.py:329" *) \$1946 ;
  assign \$1950  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1954  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h2;
  assign \$1956  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1958  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$195  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$1960  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1962  = \$1958  | (* src = "sdram_controller.py:329" *) \$1960 ;
  assign \$1964  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1968  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h2;
  assign \$1970  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1972  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1974  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1976  = \$1972  | (* src = "sdram_controller.py:329" *) \$1974 ;
  assign \$1978  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$197  = ~ (* src = "sdram_controller.py:490" *) sdramClkEn;
  assign \$1982  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h3;
  assign \$1984  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$1986  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$1988  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$1990  = \$1986  | (* src = "sdram_controller.py:329" *) \$1988 ;
  assign \$1992  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$1996  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h3;
  assign \$1998  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$1  = bankController0_bankState != (* src = "sdram_controller.py:659" *) 1'h1;
  assign \$19  = ~ (* src = "sdram_controller.py:805" *) ctrlReady;
  assign \$199  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$2000  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$2002  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$2004  = \$2000  | (* src = "sdram_controller.py:329" *) \$2002 ;
  assign \$2006  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$2010  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h3;
  assign \$2012  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$2014  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$2016  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$2018  = \$2014  | (* src = "sdram_controller.py:329" *) \$2016 ;
  assign \$201  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$2020  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$2024  = targetBankAddress == (* src = "sdram_controller.py:338" *) 2'h3;
  assign \$2026  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$2028  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$2030  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$2032  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$2034  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$2036  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$2038  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$203  = ~ (* src = "sdram_controller.py:550" *) sdramClkEn;
  assign \$2040  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$2042  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$2044  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$2046  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$2048  = \$2044  & (* src = "sdram_controller.py:613" *) \$2046 ;
  assign \$2052  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$2054  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$2056  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$2058  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$2060  = \$2056  & (* src = "sdram_controller.py:399" *) \$2058 ;
  assign \$2064  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$2066  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$2068  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$2070  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$2072  = \$2068  & (* src = "sdram_controller.py:613" *) \$2070 ;
  assign \$2076  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$2078  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$207  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$2080  = pageColumnIndex < (* src = "sdram_controller.py:913" *) 8'hff;
  assign \$2083  = pageColumnIndex + (* src = "sdram_controller.py:914" *) 1'h1;
  assign \$2085  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$2087  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$2089  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$2091  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$2094  = pageColumnIndex + (* src = "sdram_controller.py:1055" *) 1'h1;
  assign \$2096  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$2098  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$209  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$2100  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$2102  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$2104  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$2106  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$2108  = pageColumnIndex == (* src = "sdram_controller.py:1063" *) 8'hfc;
  assign \$2110  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$2112  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$2114  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$2116  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$2118  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$211  = ~ (* src = "sdram_controller.py:509" *) sdramClkEn;
  assign \$2120  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$2122  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$2124  = + (* src = "sdram_controller.py:217" *) ctrlWrDataIn;
  assign \$2126  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$2128  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$2130  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$2132  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$2134  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$2138  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$213  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$2140  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$2142  = \$2140  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  always @(posedge 1'h0)
    targetBankCanActivate <= \targetBankCanActivate$next ;
  always @(posedge 1'h0)
    targetBankCanPreCharge <= \targetBankCanPreCharge$next ;
  always @(posedge 1'h0)
    targetBankRefreshCounter <= \targetBankRefreshCounter$next ;
  always @(posedge 1'h0)
    sdramCtrlr_state <= \sdramCtrlr_state$next ;
  always @(posedge 1'h0)
    previousControllerState <= \previousControllerState$next ;
  always @(posedge 1'h0)
    currentCommand <= \currentCommand$next ;
  always @(posedge 1'h0)
    sdramClkEn <= \sdramClkEn$next ;
  always @(posedge 1'h0)
    sdramCSn <= \sdramCSn$next ;
  always @(posedge 1'h0)
    repeatRefresh <= \repeatRefresh$next ;
  always @(posedge 1'h0)
    powerUpCounter <= \powerUpCounter$next ;
  always @(posedge 1'h0)
    cmdIndex <= \cmdIndex$next ;
  always @(posedge 1'h0)
    sdramRASn <= \sdramRASn$next ;
  always @(posedge 1'h0)
    sdramCASn <= \sdramCASn$next ;
  always @(posedge 1'h0)
    sdramWEn <= \sdramWEn$next ;
  always @(posedge 1'h0)
    delayCounter <= \delayCounter$next ;
  always @(posedge 1'h0)
    sdramAddress <= \sdramAddress$next ;
  assign \$215  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  always @(posedge 1'h0)
    bankController0_bankState <= \bankController0_bankState$next ;
  always @(posedge 1'h0)
    bankController1_bankState <= \bankController1_bankState$next ;
  always @(posedge 1'h0)
    bankController2_bankState <= \bankController2_bankState$next ;
  always @(posedge 1'h0)
    bankController3_bankState <= \bankController3_bankState$next ;
  always @(posedge 1'h0)
    errorState <= \errorState$next ;
  always @(posedge 1'h0)
    sdramBank <= \sdramBank$next ;
  always @(posedge 1'h0)
    burstWritesMode <= \burstWritesMode$next ;
  always @(posedge 1'h0)
    ctrlReady <= \ctrlReady$next ;
  always @(posedge 1'h0)
    ctrlAddress <= \ctrlAddress$next ;
  always @(posedge 1'h0)
    refreshRequired <= \refreshRequired$next ;
  always @(posedge 1'h0)
    ctrlRdInProgress <= \ctrlRdInProgress$next ;
  always @(posedge 1'h0)
    sdramDataMasks <= \sdramDataMasks$next ;
  always @(posedge 1'h0)
    pageColumnIndex <= \pageColumnIndex$next ;
  always @(posedge 1'h0)
    ctrlRdIncAddress <= \ctrlRdIncAddress$next ;
  always @(posedge 1'h0)
    ctrlWrIncAddress <= \ctrlWrIncAddress$next ;
  always @(posedge 1'h0)
    sdramDqWRn <= \sdramDqWRn$next ;
  always @(posedge 1'h0)
    sdramDqIn <= \sdramDqIn$next ;
  always @(posedge 1'h0)
    ctrlWrInProgress <= \ctrlWrInProgress$next ;
  always @(posedge 1'h0)
    refreshCmdIndex <= \refreshCmdIndex$next ;
  assign \$217  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$21  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$219  = \$215  | (* src = "sdram_controller.py:329" *) \$217 ;
  assign \$221  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$225  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$227  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$229  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$231  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$233  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$235  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$237  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$23  = cmdIndex == (* src = "sdram_controller.py:935" *) 4'ha;
  assign \$239  = \$235  & (* src = "sdram_controller.py:443" *) \$237 ;
  assign \$241  = ~ (* src = "sdram_controller.py:447" *) sdramClkEn;
  assign \$243  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$245  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$247  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$249  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$251  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$253  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$255  = \$251  & (* src = "sdram_controller.py:613" *) \$253 ;
  assign \$257  = ~ (* src = "sdram_controller.py:617" *) sdramClkEn;
  assign \$25  = ! (* src = "sdram_controller.py:939" *) $signed(delayCounter);
  assign \$259  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$261  = ~ (* src = "sdram_controller.py:356" *) sdramClkEn;
  assign \$263  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$265  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$267  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$269  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$271  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$273  = \$269  | (* src = "sdram_controller.py:329" *) \$271 ;
  assign \$275  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$27  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$279  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$281  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$283  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$285  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$287  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$289  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$291  = \$287  & (* src = "sdram_controller.py:399" *) \$289 ;
  assign \$293  = ~ (* src = "sdram_controller.py:403" *) sdramClkEn;
  assign \$295  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$297  = pageColumnIndex == (* src = "sdram_controller.py:1022" *) targetColumnAddress;
  assign \$29  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$299  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$301  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$303  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$305  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$307  = \$303  & (* src = "sdram_controller.py:613" *) \$305 ;
  assign \$309  = ~ (* src = "sdram_controller.py:617" *) sdramClkEn;
  assign \$311  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$313  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$315  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$317  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$31  = ! (* src = "sdram_controller.py:1084" *) $signed(delayCounter);
  assign \$319  = ~ (* src = "sdram_controller.py:356" *) sdramClkEn;
  assign \$321  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$323  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$325  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$327  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$329  = ~ (* src = "sdram_controller.py:550" *) sdramClkEn;
  assign \$335  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$337  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$339  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$343  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$345  = ~ (* src = "sdram_controller.py:375" *) sdramClkEn;
  assign \$349  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$351  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$355  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$357  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$35  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$359  = ~ (* src = "sdram_controller.py:490" *) sdramClkEn;
  assign \$363  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$365  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$367  = ~ (* src = "sdram_controller.py:550" *) sdramClkEn;
  assign \$371  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$373  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$377  = ~ (* src = "sdram_controller.py:509" *) sdramClkEn;
  assign \$37  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$381  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$383  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$385  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$387  = \$383  | (* src = "sdram_controller.py:329" *) \$385 ;
  assign \$389  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$393  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$395  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$3  = bankController1_bankState != (* src = "sdram_controller.py:659" *) 1'h1;
  assign \$39  = \$37  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$399  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$401  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$403  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$405  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$407  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$409  = \$405  & (* src = "sdram_controller.py:443" *) \$407 ;
  assign \$411  = ~ (* src = "sdram_controller.py:447" *) sdramClkEn;
  assign \$415  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$417  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$41  = previousControllerState == (* src = "sdram_controller.py:1112" *) 3'h4;
  assign \$421  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$423  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$425  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$427  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$429  = \$425  & (* src = "sdram_controller.py:613" *) \$427 ;
  assign \$431  = ~ (* src = "sdram_controller.py:617" *) sdramClkEn;
  assign \$435  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$437  = ~ (* src = "sdram_controller.py:356" *) sdramClkEn;
  assign \$43  = previousControllerState == (* src = "sdram_controller.py:1114" *) 3'h6;
  assign \$441  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$443  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$447  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$449  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$451  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$453  = \$449  | (* src = "sdram_controller.py:329" *) \$451 ;
  assign \$455  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$45  = cmdIndex == (* src = "sdram_controller.py:726" *) 1'h1;
  assign \$459  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$461  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$465  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$467  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$469  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$471  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$473  = \$469  & (* src = "sdram_controller.py:399" *) \$471 ;
  assign \$475  = ~ (* src = "sdram_controller.py:403" *) sdramClkEn;
  assign \$47  = powerUpCounter > (* src = "sdram_controller.py:727" *) 1'h0;
  assign \$479  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$481  = pageColumnIndex == (* src = "sdram_controller.py:1022" *) targetColumnAddress;
  assign \$483  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$487  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$489  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$491  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$493  = \$489  & (* src = "sdram_controller.py:613" *) \$491 ;
  assign \$495  = ~ (* src = "sdram_controller.py:617" *) sdramClkEn;
  assign \$49  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$499  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$501  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$505  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$507  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$509  = ~ (* src = "sdram_controller.py:356" *) sdramClkEn;
  assign \$513  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$515  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$51  = ctrlWr & (* src = "sdram_controller.py:801" *) burstWritesMode;
  assign \$519  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$521  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$523  = ~ (* src = "sdram_controller.py:550" *) sdramClkEn;
  assign \$529  = ~ (* src = "sdram_controller.py:537" *) sdramClkEn;
  assign \$533  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$537  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$53  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$539  = $signed(delayCounter) > (* src = "sdram_controller.py:390" *) $signed(5'h00);
  assign \$541  = ! (* src = "sdram_controller.py:392" *) $signed(delayCounter);
  assign \$543  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$547  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$549  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$551  = $signed(delayCounter) > (* src = "sdram_controller.py:501" *) $signed(5'h00);
  assign \$553  = ! (* src = "sdram_controller.py:503" *) $signed(delayCounter);
  assign \$555  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$557  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$55  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$561  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$567  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$569  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$571  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$573  = \$569  | (* src = "sdram_controller.py:329" *) \$571 ;
  assign \$575  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$579  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$583  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$585  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$587  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$589  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$591  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$593  = \$589  & (* src = "sdram_controller.py:443" *) \$591 ;
  assign \$597  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$5  = bankController2_bankState != (* src = "sdram_controller.py:659" *) 1'h1;
  assign \$59  = $signed(delayCounter) > (* src = "sdram_controller.py:1103" *) $signed(5'h00);
  assign \$601  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$603  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$605  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$607  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$609  = \$605  & (* src = "sdram_controller.py:613" *) \$607 ;
  assign \$613  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$617  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$61  = ! (* src = "sdram_controller.py:1105" *) $signed(delayCounter);
  assign \$621  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$623  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$625  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$627  = \$623  | (* src = "sdram_controller.py:329" *) \$625 ;
  assign \$629  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$633  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$637  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$63  = \$61  & (* src = "sdram_controller.py:1105" *) cmdCompleted;
  assign \$639  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$641  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$643  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$645  = \$641  & (* src = "sdram_controller.py:399" *) \$643 ;
  assign \$649  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$651  = pageColumnIndex == (* src = "sdram_controller.py:1022" *) targetColumnAddress;
  assign \$655  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$657  = targetBankState != (* src = "sdram_controller.py:613" *) 2'h2;
  assign \$65  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$659  = targetBankState != (* src = "sdram_controller.py:614" *) 2'h3;
  assign \$661  = \$657  & (* src = "sdram_controller.py:613" *) \$659 ;
  assign \$665  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$669  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$671  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$675  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$67  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$679  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$681  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$689  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$693  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$697  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$69  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$701  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$703  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$707  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$709  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$713  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$71  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$719  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$721  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$723  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$725  = \$721  | (* src = "sdram_controller.py:329" *) \$723 ;
  assign \$727  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$731  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$735  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$737  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$73  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$739  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$741  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$743  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$745  = \$741  & (* src = "sdram_controller.py:443" *) \$743 ;
  assign \$749  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$753  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$757  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$75  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$761  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$763  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$765  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$767  = \$763  | (* src = "sdram_controller.py:329" *) \$765 ;
  assign \$769  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$773  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$777  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$77  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$779  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$781  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$783  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$785  = \$781  & (* src = "sdram_controller.py:399" *) \$783 ;
  assign \$789  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$791  = pageColumnIndex == (* src = "sdram_controller.py:1022" *) targetColumnAddress;
  assign \$795  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$7  = bankController3_bankState != (* src = "sdram_controller.py:659" *) 1'h1;
  assign \$79  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$799  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$801  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$805  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$809  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$811  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$81  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$819  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$821  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$823  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$825  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$827  = cmdIndex == (* src = "sdram_controller.py:726" *) 1'h1;
  assign \$829  = powerUpCounter > (* src = "sdram_controller.py:727" *) 1'h0;
  assign \$832  = powerUpCounter - (* src = "sdram_controller.py:728" *) 1'h1;
  assign \$834  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$836  = cmdIndex == (* src = "sdram_controller.py:726" *) 1'h1;
  assign \$838  = powerUpCounter > (* src = "sdram_controller.py:727" *) 1'h0;
  assign \$83  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$840  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$842  = cmdIndex == (* src = "sdram_controller.py:746" *) 1'h1;
  assign \$844  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$846  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$848  = cmdIndex == (* src = "sdram_controller.py:762" *) 3'h4;
  assign \$850  = cmdIndex == (* src = "sdram_controller.py:767" *) 3'h5;
  assign \$852  = $signed(delayCounter) > (* src = "sdram_controller.py:768" *) $signed(5'h00);
  assign \$854  = ! (* src = "sdram_controller.py:770" *) $signed(delayCounter);
  assign \$856  = cmdIndex == (* src = "sdram_controller.py:773" *) 3'h6;
  assign \$858  = ! (* src = "sdram_controller.py:818" *) cmdIndex;
  assign \$85  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$860  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$862  = cmdIndex == (* src = "sdram_controller.py:834" *) 2'h2;
  assign \$864  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$866  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$868  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$870  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$872  = cmdIndex == (* src = "sdram_controller.py:858" *) 3'h5;
  assign \$874  = cmdIndex == (* src = "sdram_controller.py:866" *) 3'h6;
  assign \$876  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$878  = pageColumnIndex < (* src = "sdram_controller.py:913" *) 8'hff;
  assign \$87  = cmdIndex == (* src = "sdram_controller.py:853" *) 3'h4;
  assign \$880  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$882  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$884  = cmdIndex == (* src = "sdram_controller.py:935" *) 4'ha;
  assign \$886  = ! (* src = "sdram_controller.py:939" *) $signed(delayCounter);
  assign \$888  = ! (* src = "sdram_controller.py:954" *) cmdIndex;
  assign \$890  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$892  = cmdIndex == (* src = "sdram_controller.py:967" *) 2'h2;
  assign \$894  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$896  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$898  = cmdIndex == (* src = "sdram_controller.py:1015" *) 3'h4;
  assign \$89  = cmdIndex == (* src = "sdram_controller.py:872" *) 3'h7;
  assign \$900  = pageColumnIndex < (* src = "sdram_controller.py:1054" *) 8'hff;
  assign \$902  = cmdIndex == (* src = "sdram_controller.py:1065" *) 3'h5;
  assign \$904  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$906  = cmdIndex == (* src = "sdram_controller.py:1080" *) 3'h7;
  assign \$908  = ! (* src = "sdram_controller.py:1084" *) $signed(delayCounter);
  assign \$910  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$912  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  assign \$916  = cmdIndex == (* src = "sdram_controller.py:750" *) 2'h2;
  assign \$918  = ~ (* src = "sdram_controller.py:487" *) allBanksIdle;
  assign \$91  = pageColumnIndex == (* src = "sdram_controller.py:918" *) 8'hfe;
  assign \$922  = cmdIndex == (* src = "sdram_controller.py:758" *) 2'h3;
  assign \$924  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$930  = cmdIndex == (* src = "sdram_controller.py:824" *) 1'h1;
  assign \$932  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$934  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$936  = \$932  | (* src = "sdram_controller.py:329" *) \$934 ;
  assign \$938  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$93  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$942  = cmdIndex == (* src = "sdram_controller.py:840" *) 2'h3;
  assign \$944  = $signed(delayCounter) > (* src = "sdram_controller.py:841" *) $signed(5'h00);
  assign \$946  = ! (* src = "sdram_controller.py:843" *) $signed(delayCounter);
  assign \$948  = targetBankState != (* src = "sdram_controller.py:443" *) 2'h2;
  assign \$950  = targetBankState != (* src = "sdram_controller.py:444" *) 2'h3;
  assign \$952  = \$948  & (* src = "sdram_controller.py:443" *) \$950 ;
  assign \$956  = cmdIndex == (* src = "sdram_controller.py:920" *) 4'h8;
  assign \$95  = cmdIndex == (* src = "sdram_controller.py:929" *) 4'h9;
  assign \$960  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$962  = targetBankState != (* src = "sdram_controller.py:329" *) 1'h1;
  assign \$964  = ~ (* src = "sdram_controller.py:329" *) targetBankCanActivate;
  assign \$966  = \$962  | (* src = "sdram_controller.py:329" *) \$964 ;
  assign \$968  = ~ (* src = "sdram_controller.py:331" *) sdramClkEn;
  assign \$972  = cmdIndex == (* src = "sdram_controller.py:973" *) 2'h3;
  assign \$974  = ! (* src = "sdram_controller.py:1002" *) $signed(delayCounter);
  assign \$976  = targetBankState != (* src = "sdram_controller.py:399" *) 2'h2;
  assign \$978  = targetBankState != (* src = "sdram_controller.py:400" *) 2'h3;
  assign \$97  = cmdIndex == (* src = "sdram_controller.py:958" *) 1'h1;
  assign \$980  = \$976  & (* src = "sdram_controller.py:399" *) \$978 ;
  assign \$984  = cmdIndex == (* src = "sdram_controller.py:1071" *) 3'h6;
  assign \$986  = ! (* src = "sdram_controller.py:1074" *) $signed(delayCounter);
  assign \$990  = ~ (* src = "sdram_controller.py:1096" *) refreshCmdIndex;
  assign \$992  = ~ (* src = "sdram_controller.py:547" *) allBanksIdle;
  assign \$996  = ! (* src = "sdram_controller.py:716" *) cmdIndex;
  assign \$998  = ! (* src = "sdram_controller.py:741" *) cmdIndex;
  bankController0 bankController0 (
    .bankActivated(bankController0_bankActivated),
    .bankCanActivate(bankController0_bankCanActivate),
    .bankCanPreCharge(bankController0_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController0_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController0_bankShouldRefresh),
    .bankState(bankController0_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController0_otherBankActivated)
  );
  bankController1 bankController1 (
    .bankActivated(bankController1_bankActivated),
    .bankCanActivate(bankController1_bankCanActivate),
    .bankCanPreCharge(bankController1_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController1_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController1_bankShouldRefresh),
    .bankState(bankController1_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController1_otherBankActivated)
  );
  bankController2 bankController2 (
    .bankActivated(bankController2_bankActivated),
    .bankCanActivate(bankController2_bankCanActivate),
    .bankCanPreCharge(bankController2_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController2_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController2_bankShouldRefresh),
    .bankState(bankController2_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController2_otherBankActivated)
  );
  bankController3 bankController3 (
    .bankActivated(bankController3_bankActivated),
    .bankCanActivate(bankController3_bankCanActivate),
    .bankCanPreCharge(bankController3_bankCanPreCharge),
    .bankREFIcyclesCounter(bankController3_bankREFIcyclesCounter),
    .bankShouldRefresh(bankController3_bankShouldRefresh),
    .bankState(bankController3_bankState),
    .clkSDRAM_clk(1'h0),
    .clkSDRAM_rst(1'h0),
    .otherBankActivated(bankController3_otherBankActivated)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    allBanksIdle = 1'h1;
    (* src = "sdram_controller.py:659" *)
    casez (\$1 )
      /* src = "sdram_controller.py:659" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
    (* src = "sdram_controller.py:659" *)
    casez (\$3 )
      /* src = "sdram_controller.py:659" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
    (* src = "sdram_controller.py:659" *)
    casez (\$5 )
      /* src = "sdram_controller.py:659" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
    (* src = "sdram_controller.py:659" *)
    casez (\$7 )
      /* src = "sdram_controller.py:659" */
      1'h1:
          allBanksIdle = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramCtrlr_state$next  = sdramCtrlr_state;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
        begin
          \sdramCtrlr_state$next  = 3'h0;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:726" *)
                casez (\$9 )
                  /* src = "sdram_controller.py:726" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:727" *)
                      casez (\$11 )
                        /* src = "sdram_controller.py:727" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:729" */
                        default:
                            \sdramCtrlr_state$next  = 3'h2;
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
        begin
          \sdramCtrlr_state$next  = 3'h2;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:740" */
            default:
                (* src = "sdram_controller.py:773" *)
                casez (\$13 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:776" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:776" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:779" */
                        default:
                            \sdramCtrlr_state$next  = 3'h3;
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
        begin
          \sdramCtrlr_state$next  = 3'h3;
          (* src = "sdram_controller.py:788" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:788" */
            2'b?1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:791" */
            2'b1?:
                (* src = "sdram_controller.py:792" *)
                casez ({ \$15 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:792" */
                  3'b??1:
                      \sdramCtrlr_state$next  = 3'h4;
                  /* src = "sdram_controller.py:795" */
                  3'b?1?:
                      (* src = "sdram_controller.py:799" *)
                      casez (\$17 )
                        /* src = "sdram_controller.py:799" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h5;
                      endcase
                  /* src = "sdram_controller.py:801" */
                  3'b1??:
                      (* src = "sdram_controller.py:805" *)
                      casez (\$19 )
                        /* src = "sdram_controller.py:805" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h6;
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
        begin
          \sdramCtrlr_state$next  = 3'h5;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$21 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            \sdramCtrlr_state$next  = 3'h4;
                      endcase
                endcase
                (* src = "sdram_controller.py:935" *)
                casez (\$23 )
                  /* src = "sdram_controller.py:935" */
                  1'h1:
                      (* src = "sdram_controller.py:939" *)
                      casez (\$25 )
                        /* src = "sdram_controller.py:939" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h3;
                      endcase
                endcase
              end
          endcase
        end
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
        begin
          \sdramCtrlr_state$next  = 3'h6;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$27 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            \sdramCtrlr_state$next  = 3'h4;
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$29 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      (* src = "sdram_controller.py:1084" *)
                      casez (\$31 )
                        /* src = "sdram_controller.py:1084" */
                        1'h1:
                            \sdramCtrlr_state$next  = 3'h3;
                      endcase
                endcase
              end
          endcase
        end
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
        begin
          \sdramCtrlr_state$next  = 3'h4;
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                \sdramCtrlr_state$next  = 3'h1;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1101" *)
                casez (\$33 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$39 , \$35  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:1114" *)
                            casez (\$43 )
                              /* src = "sdram_controller.py:1114" */
                              1'h1:
                                  \sdramCtrlr_state$next  = 3'h5;
                              /* src = "sdram_controller.py:1116" */
                              default:
                                  \sdramCtrlr_state$next  = 3'h3;
                            endcase
                      endcase
                endcase
          endcase
        end
      /* \amaranth.decoding  = "Error/1" */
      /* src = "sdram_controller.py:1118" */
      3'h1:
          \sdramCtrlr_state$next  = 3'h1;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramCtrlr_state$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    currentControllerState = 3'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          currentControllerState = 3'h0;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          currentControllerState = 3'h1;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          currentControllerState = 3'h2;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          currentControllerState = 3'h6;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          currentControllerState = 3'h4;
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          currentControllerState = 3'h3;
      /* \amaranth.decoding  = "Error/1" */
      /* src = "sdram_controller.py:1118" */
      3'h1:
          currentControllerState = 3'h7;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \previousControllerState$next  = previousControllerState;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:726" *)
                casez (\$45 )
                  /* src = "sdram_controller.py:726" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:727" *)
                      casez (\$47 )
                        /* src = "sdram_controller.py:727" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:729" */
                        default:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:740" */
            default:
                (* src = "sdram_controller.py:773" *)
                casez (\$49 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:776" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:776" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:779" */
                        default:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:788" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:788" */
            2'b?1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:791" */
            2'b1?:
                (* src = "sdram_controller.py:792" *)
                casez ({ \$51 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:792" */
                  3'b??1:
                      \previousControllerState$next  = currentControllerState;
                  /* src = "sdram_controller.py:795" */
                  3'b?1?:
                      \previousControllerState$next  = currentControllerState;
                  /* src = "sdram_controller.py:801" */
                  3'b1??:
                      \previousControllerState$next  = currentControllerState;
                endcase
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$53 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$55 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                \previousControllerState$next  = currentControllerState;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1101" *)
                casez (\$57 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$63 , \$59  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \previousControllerState$next  = currentControllerState;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \previousControllerState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    nextCommand = 5'h00;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$65 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$67 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      nextCommand = 5'h03;
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$69 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$71 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      nextCommand = 5'h08;
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$73 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      nextCommand = 5'h0c;
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$75 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          nextCommand = 5'h09;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$77 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            nextCommand = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$79 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$81 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$85 , \$83  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            nextCommand = 5'h06;
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$87 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$89 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$91 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            nextCommand = 5'h12;
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$93 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            nextCommand = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$95 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$97 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            nextCommand = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$99 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$101 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$103 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            nextCommand = 5'h04;
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$105 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1022" *)
                      casez (\$107 )
                        /* src = "sdram_controller.py:1022" */
                        1'h1:
                            nextCommand = 5'h0b;
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$109 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            nextCommand = 5'h12;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$111 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$113 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$115 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  nextCommand = 5'h02;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$117 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$119 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      nextCommand = 5'h0c;
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$121 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      nextCommand = 5'h0b;
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \currentCommand$next  = currentCommand;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$123 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$125 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      \currentCommand$next  = 5'h03;
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$127 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$129 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      \currentCommand$next  = 5'h08;
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$131 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      \currentCommand$next  = 5'h0c;
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$133 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          \currentCommand$next  = 5'h09;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$135 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            \currentCommand$next  = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$137 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$139 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$143 , \$141  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            \currentCommand$next  = 5'h06;
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$145 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$147 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$149 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            \currentCommand$next  = 5'h12;
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$151 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            \currentCommand$next  = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$153 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$155 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            \currentCommand$next  = 5'h01;
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$157 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$159 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$161 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            \currentCommand$next  = 5'h04;
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$163 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1022" *)
                      casez (\$165 )
                        /* src = "sdram_controller.py:1022" */
                        1'h1:
                            \currentCommand$next  = 5'h0b;
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$167 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            \currentCommand$next  = 5'h12;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$169 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$171 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$173 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  \currentCommand$next  = 5'h02;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$175 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$177 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      \currentCommand$next  = 5'h0c;
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$179 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      \currentCommand$next  = 5'h0b;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \currentCommand$next  = 5'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramClkEn$next  = sdramClkEn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$181 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$183 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \sdramClkEn$next  = 1'h0;
                      endcase
                    end
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$185 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:375" *)
                      casez (\$187 )
                        /* src = "sdram_controller.py:375" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$189 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$191 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$193 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$195 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                            (* src = "sdram_controller.py:490" *)
                            casez (\$197 )
                              /* src = "sdram_controller.py:490" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$199 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$201 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                          begin
                            (* src = "sdram_controller.py:550" *)
                            casez (\$203 )
                              /* src = "sdram_controller.py:550" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                            (* src = "sdram_controller.py:553" *)
                            casez (\$205 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$207 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$209 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:509" *)
          casez (\$211 )
            /* src = "sdram_controller.py:509" */
            1'h1:
                \sdramClkEn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$213 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$223 , \$221 , \$219  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$225 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$227 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$229 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$233 , \$231  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$239 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:447" *)
                                  casez (\$241 )
                                    /* src = "sdram_controller.py:447" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$243 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$245 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$247 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$249 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$255 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                  (* src = "sdram_controller.py:617" *)
                                  casez (\$257 )
                                    /* src = "sdram_controller.py:617" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$259 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:356" *)
                            casez (\$261 )
                              /* src = "sdram_controller.py:356" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$263 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$265 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$267 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$277 , \$275 , \$273  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$279 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$281 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$283 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$285 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$291 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:403" *)
                                  casez (\$293 )
                                    /* src = "sdram_controller.py:403" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$295 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1022" *)
                      casez (\$297 )
                        /* src = "sdram_controller.py:1022" */
                        1'h1:
                            (* src = "sdram_controller.py:537" *)
                            casez (\$299 )
                              /* src = "sdram_controller.py:537" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$301 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$307 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                  (* src = "sdram_controller.py:617" *)
                                  casez (\$309 )
                                    /* src = "sdram_controller.py:617" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$311 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$313 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$315 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$317 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:356" *)
                                  casez (\$319 )
                                    /* src = "sdram_controller.py:356" */
                                    1'h1:
                                        \sdramClkEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$321 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$323 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$325 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$327 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                          begin
                            (* src = "sdram_controller.py:550" *)
                            casez (\$329 )
                              /* src = "sdram_controller.py:550" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                            (* src = "sdram_controller.py:553" *)
                            casez (\$331 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramClkEn$next  = 1'h1;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$333 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:537" *)
                      casez (\$335 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            \sdramClkEn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramClkEn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    cmdRemainingCyclesCounter = 2'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$337 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$339 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$341 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$343 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:375" *)
                      casez (\$345 )
                        /* src = "sdram_controller.py:375" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:378" *)
                      casez (\$347 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$349 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$351 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$353 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$355 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$357 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                          begin
                            (* src = "sdram_controller.py:490" *)
                            casez (\$359 )
                              /* src = "sdram_controller.py:490" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:493" *)
                            casez (\$361 )
                              /* src = "sdram_controller.py:493" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$363 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$365 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                          begin
                            (* src = "sdram_controller.py:550" *)
                            casez (\$367 )
                              /* src = "sdram_controller.py:550" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:553" *)
                            casez (\$369 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$371 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$373 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$375 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
        begin
          (* src = "sdram_controller.py:509" *)
          casez (\$377 )
            /* src = "sdram_controller.py:509" */
            1'h1:
                cmdRemainingCyclesCounter = 2'h1;
          endcase
          (* src = "sdram_controller.py:512" *)
          casez (\$379 )
            /* src = "sdram_controller.py:512" */
            1'h1:
                cmdRemainingCyclesCounter = 2'h0;
          endcase
        end
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$381 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$391 , \$389 , \$387  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  cmdRemainingCyclesCounter = 2'h1;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$393 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$395 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$397 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$399 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$403 , \$401  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$409 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:447" *)
                                  casez (\$411 )
                                    /* src = "sdram_controller.py:447" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$413 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$415 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$417 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$419 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$421 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$423 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$429 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:617" *)
                                  casez (\$431 )
                                    /* src = "sdram_controller.py:617" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:620" *)
                                  casez (\$433 )
                                    /* src = "sdram_controller.py:620" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$435 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                          begin
                            (* src = "sdram_controller.py:356" *)
                            casez (\$437 )
                              /* src = "sdram_controller.py:356" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:359" *)
                            casez (\$439 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$441 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$443 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$445 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$447 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$457 , \$455 , \$453  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  cmdRemainingCyclesCounter = 2'h1;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$459 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$461 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$463 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$465 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$467 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$473 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:403" *)
                                  casez (\$475 )
                                    /* src = "sdram_controller.py:403" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$477 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$479 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1022" *)
                      casez (\$481 )
                        /* src = "sdram_controller.py:1022" */
                        1'h1:
                          begin
                            (* src = "sdram_controller.py:537" *)
                            casez (\$483 )
                              /* src = "sdram_controller.py:537" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:540" *)
                            casez (\$485 )
                              /* src = "sdram_controller.py:540" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$487 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$493 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                begin
                                  (* src = "sdram_controller.py:617" *)
                                  casez (\$495 )
                                    /* src = "sdram_controller.py:617" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:620" *)
                                  casez (\$497 )
                                    /* src = "sdram_controller.py:620" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$499 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$501 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$503 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$505 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$507 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                begin
                                  (* src = "sdram_controller.py:356" *)
                                  casez (\$509 )
                                    /* src = "sdram_controller.py:356" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h1;
                                  endcase
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$511 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        cmdRemainingCyclesCounter = 2'h0;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$513 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$515 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$517 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$519 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$521 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                          begin
                            (* src = "sdram_controller.py:550" *)
                            casez (\$523 )
                              /* src = "sdram_controller.py:550" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h1;
                            endcase
                            (* src = "sdram_controller.py:553" *)
                            casez (\$525 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  cmdRemainingCyclesCounter = 2'h0;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$527 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:537" *)
                      casez (\$529 )
                        /* src = "sdram_controller.py:537" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h1;
                      endcase
                      (* src = "sdram_controller.py:540" *)
                      casez (\$531 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdRemainingCyclesCounter = 2'h0;
                      endcase
                    end
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    cmdCompleted = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$533 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$535 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$537 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:390" *)
                      casez ({ \$541 , \$539  })
                        /* src = "sdram_controller.py:390" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:392" */
                        2'b1?:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$543 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$545 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$547 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$549 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                            (* src = "sdram_controller.py:501" *)
                            casez ({ \$553 , \$551  })
                              /* src = "sdram_controller.py:501" */
                              2'b?1:
                                  /* empty */;
                              /* src = "sdram_controller.py:503" */
                              2'b1?:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$555 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$557 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$559 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$561 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$563 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:512" *)
          casez (\$565 )
            /* src = "sdram_controller.py:512" */
            1'h1:
                cmdCompleted = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$567 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$577 , \$575 , \$573  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$579 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$581 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$583 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$587 , \$585  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$593 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$595 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$597 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$599 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$601 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$603 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$609 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                  (* src = "sdram_controller.py:620" *)
                                  casez (\$611 )
                                    /* src = "sdram_controller.py:620" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$613 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$615 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$617 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$619 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$621 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$631 , \$629 , \$627  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$633 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$635 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$637 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$639 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$645 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$647 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$649 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1022" *)
                      casez (\$651 )
                        /* src = "sdram_controller.py:1022" */
                        1'h1:
                            (* src = "sdram_controller.py:540" *)
                            casez (\$653 )
                              /* src = "sdram_controller.py:540" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$655 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$661 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                  (* src = "sdram_controller.py:620" *)
                                  casez (\$663 )
                                    /* src = "sdram_controller.py:620" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$665 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$667 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$669 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$671 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$673 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        cmdCompleted = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$675 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$677 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$679 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$681 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$683 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  cmdCompleted = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$685 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$687 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            cmdCompleted = 1'h1;
                      endcase
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramCSn$next  = sdramCSn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$689 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$691 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$693 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$695 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \sdramCSn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$697 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$699 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$701 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$703 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                            (* src = "sdram_controller.py:493" *)
                            casez (\$705 )
                              /* src = "sdram_controller.py:493" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$707 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$709 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$711 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$713 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$715 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:512" *)
          casez (\$717 )
            /* src = "sdram_controller.py:512" */
            1'h1:
                \sdramCSn$next  = 1'h0;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$719 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$729 , \$727 , \$725  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$731 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$733 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$735 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$739 , \$737  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$745 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$747 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        \sdramCSn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$749 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$751 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$753 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$755 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$757 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$759 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$761 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$771 , \$769 , \$767  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$773 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$775 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$777 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$779 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$785 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$787 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramCSn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$789 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* src = "sdram_controller.py:1022" *)
                      casez (\$791 )
                        /* src = "sdram_controller.py:1022" */
                        1'h1:
                            (* src = "sdram_controller.py:540" *)
                            casez (\$793 )
                              /* src = "sdram_controller.py:540" */
                              1'h1:
                                  \sdramCSn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$795 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$797 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$799 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$801 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$803 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \sdramCSn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$805 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$807 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$809 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$811 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$813 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramCSn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$815 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:540" *)
                      casez (\$817 )
                        /* src = "sdram_controller.py:540" */
                        1'h1:
                            \sdramCSn$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramCSn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    banksShouldRefresh = 1'h0;
    (* src = "sdram_controller.py:663" *)
    casez (bankController0_bankShouldRefresh)
      /* src = "sdram_controller.py:663" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
    (* src = "sdram_controller.py:663" *)
    casez (bankController1_bankShouldRefresh)
      /* src = "sdram_controller.py:663" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
    (* src = "sdram_controller.py:663" *)
    casez (bankController2_bankShouldRefresh)
      /* src = "sdram_controller.py:663" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
    (* src = "sdram_controller.py:663" *)
    casez (bankController3_bankShouldRefresh)
      /* src = "sdram_controller.py:663" */
      1'h1:
          banksShouldRefresh = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \repeatRefresh$next  = repeatRefresh;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$819 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \repeatRefresh$next  = 1'h0;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$821 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:743" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:743" */
                        1'h1:
                            \repeatRefresh$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:773" *)
                casez (\$823 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      (* src = "sdram_controller.py:776" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:776" */
                        1'h1:
                            \repeatRefresh$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \repeatRefresh$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \powerUpCounter$next  = powerUpCounter;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
              begin
                (* src = "sdram_controller.py:716" *)
                casez (\$825 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \powerUpCounter$next  = 15'h5dc0;
                      endcase
                endcase
                (* src = "sdram_controller.py:726" *)
                casez (\$827 )
                  /* src = "sdram_controller.py:726" */
                  1'h1:
                      (* src = "sdram_controller.py:727" *)
                      casez (\$829 )
                        /* src = "sdram_controller.py:727" */
                        1'h1:
                            \powerUpCounter$next  = \$832 [14:0];
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \powerUpCounter$next  = 15'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \cmdIndex$next  = cmdIndex;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
              begin
                (* src = "sdram_controller.py:716" *)
                casez (\$834 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \cmdIndex$next  = 4'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:726" *)
                casez (\$836 )
                  /* src = "sdram_controller.py:726" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:727" *)
                      casez (\$838 )
                        /* src = "sdram_controller.py:727" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:729" */
                        default:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$840 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:743" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:743" */
                        1'h1:
                            \cmdIndex$next  = 4'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:746" *)
                casez (\$842 )
                  /* src = "sdram_controller.py:746" */
                  1'h1:
                      (* src = "sdram_controller.py:748" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:748" */
                        1'h1:
                            \cmdIndex$next  = 4'h2;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$844 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* src = "sdram_controller.py:755" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:755" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$846 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:760" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:760" */
                        1'h1:
                            \cmdIndex$next  = 4'h4;
                      endcase
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$848 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      (* src = "sdram_controller.py:764" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:764" */
                        1'h1:
                            \cmdIndex$next  = 4'h5;
                      endcase
                endcase
                (* src = "sdram_controller.py:767" *)
                casez (\$850 )
                  /* src = "sdram_controller.py:767" */
                  1'h1:
                      (* src = "sdram_controller.py:768" *)
                      casez ({ \$854 , \$852  })
                        /* src = "sdram_controller.py:768" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:770" */
                        2'b1?:
                            \cmdIndex$next  = 4'h6;
                      endcase
                endcase
                (* src = "sdram_controller.py:773" *)
                casez (\$856 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:776" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:776" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                        /* src = "sdram_controller.py:779" */
                        default:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:818" *)
                casez (\$858 )
                  /* src = "sdram_controller.py:818" */
                  1'h1:
                      \cmdIndex$next  = 4'h1;
                endcase
                (* src = "sdram_controller.py:824" *)
                casez (\$860 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:832" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:832" */
                              1'h1:
                                  \cmdIndex$next  = 4'h2;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:834" *)
                casez (\$862 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      (* src = "sdram_controller.py:837" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:837" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$864 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$868 , \$866  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* src = "sdram_controller.py:849" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:849" */
                              1'h1:
                                  \cmdIndex$next  = 4'h4;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:853" *)
                casez (\$870 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      (* src = "sdram_controller.py:855" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:855" */
                        1'h1:
                            \cmdIndex$next  = 4'h5;
                      endcase
                endcase
                (* src = "sdram_controller.py:858" *)
                casez (\$872 )
                  /* src = "sdram_controller.py:858" */
                  1'h1:
                      \cmdIndex$next  = 4'h6;
                endcase
                (* src = "sdram_controller.py:866" *)
                casez (\$874 )
                  /* src = "sdram_controller.py:866" */
                  1'h1:
                      \cmdIndex$next  = 4'h7;
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$876 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:913" *)
                      casez (\$878 )
                        /* src = "sdram_controller.py:913" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:915" */
                        default:
                            \cmdIndex$next  = 4'h8;
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$880 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:927" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:927" */
                              1'h1:
                                  \cmdIndex$next  = 4'h9;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$882 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      (* src = "sdram_controller.py:932" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:932" */
                        1'h1:
                            \cmdIndex$next  = 4'ha;
                      endcase
                endcase
                (* src = "sdram_controller.py:935" *)
                casez (\$884 )
                  /* src = "sdram_controller.py:935" */
                  1'h1:
                      (* src = "sdram_controller.py:939" *)
                      casez (\$886 )
                        /* src = "sdram_controller.py:939" */
                        1'h1:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:954" *)
                casez (\$888 )
                  /* src = "sdram_controller.py:954" */
                  1'h1:
                      \cmdIndex$next  = 4'h1;
                endcase
                (* src = "sdram_controller.py:958" *)
                casez (\$890 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:965" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:965" */
                              1'h1:
                                  \cmdIndex$next  = 4'h2;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:967" *)
                casez (\$892 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      (* src = "sdram_controller.py:969" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:969" */
                        1'h1:
                            \cmdIndex$next  = 4'h3;
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$894 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$896 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* src = "sdram_controller.py:1010" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1010" */
                              1'h1:
                                  \cmdIndex$next  = 4'h4;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$898 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$900 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* src = "sdram_controller.py:1059" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1059" */
                              1'h1:
                                  \cmdIndex$next  = 4'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$902 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      (* src = "sdram_controller.py:1069" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1069" */
                        1'h1:
                            \cmdIndex$next  = 4'h6;
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$904 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1078" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1078" */
                        1'h1:
                            \cmdIndex$next  = 4'h7;
                      endcase
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$906 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      (* src = "sdram_controller.py:1084" *)
                      casez (\$908 )
                        /* src = "sdram_controller.py:1084" */
                        1'h1:
                            \cmdIndex$next  = 4'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \cmdIndex$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramRASn$next  = sdramRASn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$910 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \sdramRASn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$912 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$914 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \sdramRASn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$916 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$918 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                            (* src = "sdram_controller.py:493" *)
                            casez (\$920 )
                              /* src = "sdram_controller.py:493" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$922 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$924 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$926 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:512" *)
          casez (\$928 )
            /* src = "sdram_controller.py:512" */
            1'h1:
                \sdramRASn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$930 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$940 , \$938 , \$936  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$942 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$946 , \$944  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$952 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$954 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        \sdramRASn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$956 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$958 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$960 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$970 , \$968 , \$966  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$972 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$974 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$980 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$982 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramRASn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$984 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$986 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$988 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \sdramRASn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1096" *)
                casez (\$990 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$992 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$994 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramRASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramRASn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramCASn$next  = sdramCASn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$996 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \sdramCASn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$998 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1000 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \sdramCASn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$1002 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$1004 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                            (* src = "sdram_controller.py:493" *)
                            casez (\$1006 )
                              /* src = "sdram_controller.py:493" */
                              1'h1:
                                  \sdramCASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1008 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1010 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1012 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramCASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:512" *)
          casez (\$1014 )
            /* src = "sdram_controller.py:512" */
            1'h1:
                \sdramCASn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1016 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1026 , \$1024 , \$1022  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramCASn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$1028 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$1032 , \$1030  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$1038 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$1040 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        \sdramCASn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1042 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1044 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  \sdramCASn$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1046 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1056 , \$1054 , \$1052  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramCASn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$1058 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$1060 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$1066 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$1068 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramCASn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1070 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1072 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1074 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \sdramCASn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1096" *)
                casez (\$1076 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1078 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1080 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramCASn$next  = 1'h0;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramCASn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramWEn$next  = sdramWEn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:716" *)
                casez (\$1082 )
                  /* src = "sdram_controller.py:716" */
                  1'h1:
                      (* src = "sdram_controller.py:718" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:718" */
                        1'h1:
                            \sdramWEn$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1084 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1086 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \sdramWEn$next  = 1'h0;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$1088 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$1090 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                            (* src = "sdram_controller.py:493" *)
                            casez (\$1092 )
                              /* src = "sdram_controller.py:493" */
                              1'h1:
                                  \sdramWEn$next  = 1'h0;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1094 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1096 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1098 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:512" *)
          casez (\$1100 )
            /* src = "sdram_controller.py:512" */
            1'h1:
                \sdramWEn$next  = 1'h1;
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1102 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1112 , \$1110 , \$1108  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$1114 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$1118 , \$1116  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$1124 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$1126 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        \sdramWEn$next  = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1128 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1130 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  \sdramWEn$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1132 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1142 , \$1140 , \$1138  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$1144 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$1146 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$1152 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$1154 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramWEn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1156 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1158 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1160 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \sdramWEn$next  = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1096" *)
                casez (\$1162 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1164 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1166 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \sdramWEn$next  = 1'h1;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramWEn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \delayCounter$next  = delayCounter;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:712" *)
          casez (errorState)
            /* src = "sdram_controller.py:712" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:715" */
            default:
                (* src = "sdram_controller.py:726" *)
                casez (\$1168 )
                  /* src = "sdram_controller.py:726" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:727" *)
                      casez (\$1170 )
                        /* src = "sdram_controller.py:727" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:729" */
                        default:
                            \delayCounter$next  = 5'h1f;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1172 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1174 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \delayCounter$next  = 5'h02;
                      endcase
                      (* src = "sdram_controller.py:390" *)
                      casez ({ \$1178 , \$1176  })
                        /* src = "sdram_controller.py:390" */
                        2'b?1:
                            \delayCounter$next  = \$1181 [4:0];
                        /* src = "sdram_controller.py:392" */
                        2'b1?:
                            \delayCounter$next  = 5'h1f;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$1183 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:487" *)
                      casez (\$1185 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:489" */
                        default:
                          begin
                            (* src = "sdram_controller.py:493" *)
                            casez (\$1187 )
                              /* src = "sdram_controller.py:493" */
                              1'h1:
                                  \delayCounter$next  = 5'h01;
                            endcase
                            (* src = "sdram_controller.py:501" *)
                            casez ({ \$1191 , \$1189  })
                              /* src = "sdram_controller.py:501" */
                              2'b?1:
                                  \delayCounter$next  = \$1194 [4:0];
                              /* src = "sdram_controller.py:503" */
                              2'b1?:
                                  \delayCounter$next  = 5'h1f;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:762" *)
                casez (\$1196 )
                  /* src = "sdram_controller.py:762" */
                  1'h1:
                      (* src = "sdram_controller.py:764" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:764" */
                        1'h1:
                            \delayCounter$next  = 5'h07;
                      endcase
                endcase
                (* src = "sdram_controller.py:767" *)
                casez (\$1198 )
                  /* src = "sdram_controller.py:767" */
                  1'h1:
                      (* src = "sdram_controller.py:768" *)
                      casez ({ \$1202 , \$1200  })
                        /* src = "sdram_controller.py:768" */
                        2'b?1:
                            \delayCounter$next  = \$1205 [4:0];
                        /* src = "sdram_controller.py:770" */
                        2'b1?:
                            \delayCounter$next  = 5'h1f;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:834" *)
                casez (\$1207 )
                  /* src = "sdram_controller.py:834" */
                  1'h1:
                      (* src = "sdram_controller.py:837" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:837" */
                        1'h1:
                            \delayCounter$next  = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$1209 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$1213 , \$1211  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            \delayCounter$next  = \$1216 [4:0];
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            \delayCounter$next  = 5'h1f;
                      endcase
                endcase
                (* src = "sdram_controller.py:929" *)
                casez (\$1218 )
                  /* src = "sdram_controller.py:929" */
                  1'h1:
                      (* src = "sdram_controller.py:932" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:932" */
                        1'h1:
                            \delayCounter$next  = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:935" *)
                casez (\$1220 )
                  /* src = "sdram_controller.py:935" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:937" *)
                      casez (\$1222 )
                        /* src = "sdram_controller.py:937" */
                        1'h1:
                            \delayCounter$next  = \$1225 [4:0];
                      endcase
                      (* src = "sdram_controller.py:939" *)
                      casez (\$1227 )
                        /* src = "sdram_controller.py:939" */
                        1'h1:
                            \delayCounter$next  = 5'h1f;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:967" *)
                casez (\$1229 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      (* src = "sdram_controller.py:969" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:969" */
                        1'h1:
                            \delayCounter$next  = 5'h02;
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$1231 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1000" *)
                      casez (\$1233 )
                        /* src = "sdram_controller.py:1000" */
                        1'h1:
                            \delayCounter$next  = \$1236 [4:0];
                      endcase
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$1238 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            \delayCounter$next  = 5'h1f;
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$1240 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$1242 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* src = "sdram_controller.py:1059" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1059" */
                              1'h1:
                                  \delayCounter$next  = 5'h00;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1065" *)
                casez (\$1244 )
                  /* src = "sdram_controller.py:1065" */
                  1'h1:
                      (* src = "sdram_controller.py:1067" *)
                      casez (\$1246 )
                        /* src = "sdram_controller.py:1067" */
                        1'h1:
                            \delayCounter$next  = \$1249 [4:0];
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1251 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1072" *)
                      casez (\$1253 )
                        /* src = "sdram_controller.py:1072" */
                        1'h1:
                            \delayCounter$next  = \$1256 [4:0];
                      endcase
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1258 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  \delayCounter$next  = 5'h02;
                            endcase
                      endcase
                    end
                endcase
                (* src = "sdram_controller.py:1080" *)
                casez (\$1260 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                    begin
                      (* src = "sdram_controller.py:1082" *)
                      casez (\$1262 )
                        /* src = "sdram_controller.py:1082" */
                        1'h1:
                            \delayCounter$next  = \$1265 [4:0];
                      endcase
                      (* src = "sdram_controller.py:1084" *)
                      casez (\$1267 )
                        /* src = "sdram_controller.py:1084" */
                        1'h1:
                            \delayCounter$next  = 5'h1f;
                      endcase
                    end
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$1269 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* src = "sdram_controller.py:1098" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1098" */
                        1'h1:
                            \delayCounter$next  = 5'h07;
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$1271 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$1277 , \$1273  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            \delayCounter$next  = \$1280 [4:0];
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \delayCounter$next  = 5'h1f;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \delayCounter$next  = 5'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramAddress$next  = sdramAddress;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1282 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1284 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \sdramAddress$next [10] = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:750" *)
                casez (\$1286 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* src = "sdram_controller.py:752" *)
                      casez (\$1288 )
                        /* src = "sdram_controller.py:752" */
                        1'h1:
                          begin
                            \sdramAddress$next [10] = 1'h0;
                            \sdramAddress$next [9] = 1'h0;
                            \sdramAddress$next [8:7] = 2'h0;
                            \sdramAddress$next [6:4] = 3'h3;
                            \sdramAddress$next [3] = 1'h0;
                            \sdramAddress$next [2:0] = 3'h7;
                          end
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1290 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1300 , \$1298 , \$1296  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramAddress$next  = targetRowAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$1302 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$1306 , \$1304  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$1312 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$1314 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        \sdramAddress$next  = { 3'h0, targetColumnAddress };
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1316 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1318 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  \sdramAddress$next [10] = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1320 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1330 , \$1328 , \$1326  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramAddress$next  = targetRowAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$1332 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$1334 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$1340 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$1342 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramAddress$next  = { 3'h0, targetColumnAddress };
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1344 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1346 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1348 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        \sdramAddress$next [10] = 1'h0;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramAddress$next  = 11'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController0_bankState$next  = bankController0_bankState;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1350 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1352 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \bankController0_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1354 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1356 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1358 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController0_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:773" *)
                casez (\$1360 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      \bankController0_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1362 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1372 , \$1370 , \$1368  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1374 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController0_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController0_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1376 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1378 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  (* src = "sdram_controller.py:363" *)
                                  casez (\$1380 )
                                    /* src = "sdram_controller.py:363" */
                                    1'h1:
                                        \bankController0_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1382 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1392 , \$1390 , \$1388  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1394 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController0_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController0_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1396 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1398 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1400 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        (* src = "sdram_controller.py:363" *)
                                        casez (\$1402 )
                                          /* src = "sdram_controller.py:363" */
                                          1'h1:
                                              \bankController0_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$1404 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1406 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1408 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController0_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$1410 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$1416 , \$1412  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \bankController0_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController0_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController1_bankState$next  = bankController1_bankState;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1418 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1420 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \bankController1_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1422 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1424 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1426 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController1_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:773" *)
                casez (\$1428 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      \bankController1_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1430 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1440 , \$1438 , \$1436  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1442 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController1_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController1_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1444 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1446 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  (* src = "sdram_controller.py:363" *)
                                  casez (\$1448 )
                                    /* src = "sdram_controller.py:363" */
                                    1'h1:
                                        \bankController1_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1450 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1460 , \$1458 , \$1456  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1462 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController1_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController1_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1464 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1466 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1468 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        (* src = "sdram_controller.py:363" *)
                                        casez (\$1470 )
                                          /* src = "sdram_controller.py:363" */
                                          1'h1:
                                              \bankController1_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$1472 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1474 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1476 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController1_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$1478 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$1484 , \$1480  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \bankController1_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController1_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:667" *)
    casez (targetBankAddress)
      2'h0:
          targetBankState = bankController0_bankState;
      2'h1:
          targetBankState = bankController1_bankState;
      2'h2:
          targetBankState = bankController2_bankState;
      2'h?:
          targetBankState = bankController3_bankState;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController2_bankState$next  = bankController2_bankState;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1486 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1488 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \bankController2_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1490 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1492 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1494 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController2_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:773" *)
                casez (\$1496 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      \bankController2_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1498 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1508 , \$1506 , \$1504  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1510 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController2_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController2_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1512 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1514 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  (* src = "sdram_controller.py:363" *)
                                  casez (\$1516 )
                                    /* src = "sdram_controller.py:363" */
                                    1'h1:
                                        \bankController2_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1518 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1528 , \$1526 , \$1524  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1530 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController2_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController2_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1532 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1534 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1536 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        (* src = "sdram_controller.py:363" *)
                                        casez (\$1538 )
                                          /* src = "sdram_controller.py:363" */
                                          1'h1:
                                              \bankController2_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$1540 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1542 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1544 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController2_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$1546 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$1552 , \$1548  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \bankController2_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController2_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \bankController3_bankState$next  = bankController3_bankState;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:741" *)
                casez (\$1554 )
                  /* src = "sdram_controller.py:741" */
                  1'h1:
                      (* src = "sdram_controller.py:378" *)
                      casez (\$1556 )
                        /* src = "sdram_controller.py:378" */
                        1'h1:
                            \bankController3_bankState$next  = 3'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1558 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1560 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1562 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController3_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:773" *)
                casez (\$1564 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      \bankController3_bankState$next  = 3'h1;
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1566 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1576 , \$1574 , \$1572  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1578 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController3_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController3_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$1580 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      (* src = "sdram_controller.py:925" *)
                      casez (targetBankCanPreCharge)
                        /* src = "sdram_controller.py:925" */
                        1'h1:
                            (* src = "sdram_controller.py:359" *)
                            casez (\$1582 )
                              /* src = "sdram_controller.py:359" */
                              1'h1:
                                  (* src = "sdram_controller.py:363" *)
                                  casez (\$1584 )
                                    /* src = "sdram_controller.py:363" */
                                    1'h1:
                                        \bankController3_bankState$next  = 3'h1;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1586 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1596 , \$1594 , \$1592  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1598 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        (* full_case = 32'd1 *)
                                        (* src = "sdram_controller.py:340" *)
                                        casez (burstWritesMode)
                                          /* src = "sdram_controller.py:340" */
                                          1'h1:
                                              \bankController3_bankState$next  = 3'h3;
                                          /* src = "sdram_controller.py:342" */
                                          default:
                                              \bankController3_bankState$next  = 3'h2;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1071" *)
                casez (\$1600 )
                  /* src = "sdram_controller.py:1071" */
                  1'h1:
                      (* src = "sdram_controller.py:1074" *)
                      casez (\$1602 )
                        /* src = "sdram_controller.py:1074" */
                        1'h1:
                            (* src = "sdram_controller.py:1075" *)
                            casez (targetBankCanPreCharge)
                              /* src = "sdram_controller.py:1075" */
                              1'h1:
                                  (* src = "sdram_controller.py:359" *)
                                  casez (\$1604 )
                                    /* src = "sdram_controller.py:359" */
                                    1'h1:
                                        (* src = "sdram_controller.py:363" *)
                                        casez (\$1606 )
                                          /* src = "sdram_controller.py:363" */
                                          1'h1:
                                              \bankController3_bankState$next  = 3'h1;
                                        endcase
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$1608 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1610 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:549" */
                        default:
                            (* src = "sdram_controller.py:553" *)
                            casez (\$1612 )
                              /* src = "sdram_controller.py:553" */
                              1'h1:
                                  \bankController3_bankState$next  = 3'h5;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$1614 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$1620 , \$1616  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \bankController3_bankState$next  = 3'h1;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \bankController3_bankState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \errorState$next  = errorState;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
              begin
                (* src = "sdram_controller.py:750" *)
                casez (\$1622 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* src = "sdram_controller.py:487" *)
                      casez (\$1624 )
                        /* src = "sdram_controller.py:487" */
                        1'h1:
                            \errorState$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:758" *)
                casez (\$1626 )
                  /* src = "sdram_controller.py:758" */
                  1'h1:
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1628 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            \errorState$next  = 1'h1;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1630 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1640 , \$1638 , \$1636  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$1642 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$1646 , \$1644  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* src = "sdram_controller.py:443" *)
                            casez (\$1652 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$1654 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$1656 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            (* src = "sdram_controller.py:613" *)
                            casez (\$1662 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1664 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1674 , \$1672 , \$1670  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$1676 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$1678 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* src = "sdram_controller.py:399" *)
                            casez (\$1684 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$1686 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$1688 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* src = "sdram_controller.py:613" *)
                            casez (\$1694 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  \errorState$next  = 1'h1;
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1096" *)
                casez (\$1696 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* src = "sdram_controller.py:547" *)
                      casez (\$1698 )
                        /* src = "sdram_controller.py:547" */
                        1'h1:
                            \errorState$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \errorState$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramBank$next  = sdramBank;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
                (* src = "sdram_controller.py:750" *)
                casez (\$1700 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* src = "sdram_controller.py:752" *)
                      casez (\$1702 )
                        /* src = "sdram_controller.py:752" */
                        1'h1:
                            \sdramBank$next  = 2'h0;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:824" *)
                casez (\$1704 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1714 , \$1712 , \$1710  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramBank$next  = targetBankAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:840" *)
                casez (\$1716 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$1720 , \$1718  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:443" *)
                            casez (\$1726 )
                              /* src = "sdram_controller.py:443" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:446" */
                              default:
                                  (* src = "sdram_controller.py:450" *)
                                  casez (\$1728 )
                                    /* src = "sdram_controller.py:450" */
                                    1'h1:
                                        \sdramBank$next  = targetBankAddress;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:958" *)
                casez (\$1730 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1740 , \$1738 , \$1736  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  \sdramBank$next  = targetBankAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:973" *)
                casez (\$1742 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$1744 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$1750 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$1752 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramBank$next  = targetBankAddress;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramBank$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \burstWritesMode$next  = burstWritesMode;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
                (* src = "sdram_controller.py:750" *)
                casez (\$1754 )
                  /* src = "sdram_controller.py:750" */
                  1'h1:
                      (* src = "sdram_controller.py:755" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:755" */
                        1'h1:
                            \burstWritesMode$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \burstWritesMode$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlReady$next  = ctrlReady;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:737" *)
          casez (errorState)
            /* src = "sdram_controller.py:737" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:740" */
            default:
                (* src = "sdram_controller.py:773" *)
                casez (\$1756 )
                  /* src = "sdram_controller.py:773" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:776" *)
                      casez (repeatRefresh)
                        /* src = "sdram_controller.py:776" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:779" */
                        default:
                            \ctrlReady$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:788" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:788" */
            2'b?1:
                /* empty */;
            /* src = "sdram_controller.py:791" */
            2'b1?:
                (* src = "sdram_controller.py:792" *)
                casez ({ \$1758 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:792" */
                  3'b??1:
                      /* empty */;
                  /* src = "sdram_controller.py:795" */
                  3'b?1?:
                      \ctrlReady$next  = 1'h0;
                  /* src = "sdram_controller.py:801" */
                  3'b1??:
                      \ctrlReady$next  = 1'h0;
                endcase
          endcase
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:935" *)
                casez (\$1760 )
                  /* src = "sdram_controller.py:935" */
                  1'h1:
                      (* src = "sdram_controller.py:939" *)
                      casez (\$1762 )
                        /* src = "sdram_controller.py:939" */
                        1'h1:
                            \ctrlReady$next  = 1'h1;
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:1080" *)
                casez (\$1764 )
                  /* src = "sdram_controller.py:1080" */
                  1'h1:
                      (* src = "sdram_controller.py:1084" *)
                      casez (\$1766 )
                        /* src = "sdram_controller.py:1084" */
                        1'h1:
                            \ctrlReady$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlReady$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlAddress$next  = ctrlAddress;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          (* src = "sdram_controller.py:788" *)
          casez ({ cmdCompleted, errorState })
            /* src = "sdram_controller.py:788" */
            2'b?1:
                /* empty */;
            /* src = "sdram_controller.py:791" */
            2'b1?:
                (* src = "sdram_controller.py:792" *)
                casez ({ \$1768 , ctrlRd, banksShouldRefresh })
                  /* src = "sdram_controller.py:792" */
                  3'b??1:
                      /* empty */;
                  /* src = "sdram_controller.py:795" */
                  3'b?1?:
                      \ctrlAddress$next  = ctrlRdAddress;
                  /* src = "sdram_controller.py:801" */
                  3'b1??:
                      \ctrlAddress$next  = ctrlWrAddress;
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlAddress$next  = 21'h000000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \refreshRequired$next  = refreshRequired;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:818" *)
                casez (\$1770 )
                  /* src = "sdram_controller.py:818" */
                  1'h1:
                      \refreshRequired$next  = \$1780 ;
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:954" *)
                casez (\$1782 )
                  /* src = "sdram_controller.py:954" */
                  1'h1:
                      \refreshRequired$next  = \$1792 ;
                endcase
          endcase
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
                (* src = "sdram_controller.py:1101" *)
                casez (\$1794 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$1800 , \$1796  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \refreshRequired$next  = 1'h0;
                      endcase
                endcase
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \refreshRequired$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController0_bankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1802 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1812 , \$1810 , \$1808  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1814 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController0_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1816 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1826 , \$1824 , \$1822  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1828 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController0_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController0_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1830 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1840 , \$1838 , \$1836  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1842 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController0_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1844 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1854 , \$1852 , \$1850  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1856 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController0_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:668" *)
    casez (targetBankAddress)
      2'h0:
          \targetBankCanActivate$next  = bankController0_bankCanActivate;
      2'h1:
          \targetBankCanActivate$next  = bankController1_bankCanActivate;
      2'h2:
          \targetBankCanActivate$next  = bankController2_bankCanActivate;
      2'h?:
          \targetBankCanActivate$next  = bankController3_bankCanActivate;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \targetBankCanActivate$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController1_bankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1858 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1868 , \$1866 , \$1864  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1870 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController1_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1872 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1882 , \$1880 , \$1878  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1884 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController1_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController1_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1886 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1896 , \$1894 , \$1892  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1898 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController1_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1900 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1910 , \$1908 , \$1906  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1912 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController1_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController2_bankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1914 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1924 , \$1922 , \$1920  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1926 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController2_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1928 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1938 , \$1936 , \$1934  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1940 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController2_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController2_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1942 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1952 , \$1950 , \$1948  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1954 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController2_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1956 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1966 , \$1964 , \$1962  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1968 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController2_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController3_bankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1970 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1980 , \$1978 , \$1976  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1982 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController3_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$1984 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$1994 , \$1992 , \$1990  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$1996 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        bankController3_bankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    bankController3_otherBankActivated = 1'h0;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
                (* src = "sdram_controller.py:824" *)
                casez (\$1998 )
                  /* src = "sdram_controller.py:824" */
                  1'h1:
                      (* src = "sdram_controller.py:826" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:826" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:830" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$2008 , \$2006 , \$2004  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$2010 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController3_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
                (* src = "sdram_controller.py:958" *)
                casez (\$2012 )
                  /* src = "sdram_controller.py:958" */
                  1'h1:
                      (* src = "sdram_controller.py:959" *)
                      casez ({ targetBankCanActivate, refreshRequired })
                        /* src = "sdram_controller.py:959" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:963" */
                        2'b1?:
                            (* src = "sdram_controller.py:329" *)
                            casez ({ \$2022 , \$2020 , \$2018  })
                              /* src = "sdram_controller.py:329" */
                              3'b??1:
                                  /* empty */;
                              /* src = "sdram_controller.py:331" */
                              3'b?1?:
                                  /* empty */;
                              /* src = "sdram_controller.py:334" */
                              3'b1??:
                                  (* full_case = 32'd1 *)
                                  (* src = "sdram_controller.py:338" *)
                                  casez (\$2024 )
                                    /* src = "sdram_controller.py:338" */
                                    1'h1:
                                        /* empty */;
                                    /* src = "sdram_controller.py:344" */
                                    default:
                                        bankController3_otherBankActivated = 1'h1;
                                  endcase
                            endcase
                      endcase
                endcase
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlRdInProgress$next  = ctrlRdInProgress;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:840" *)
                casez (\$2026 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$2030 , \$2028  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* src = "sdram_controller.py:849" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:849" */
                              1'h1:
                                  \ctrlRdInProgress$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$2032 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      \ctrlRdInProgress$next  = 1'h0;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlRdInProgress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramDataMasks$next  = sdramDataMasks;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:840" *)
                casez (\$2034 )
                  /* src = "sdram_controller.py:840" */
                  1'h1:
                      (* src = "sdram_controller.py:841" *)
                      casez ({ \$2038 , \$2036  })
                        /* src = "sdram_controller.py:841" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:843" */
                        2'b1?:
                            (* src = "sdram_controller.py:849" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:849" */
                              1'h1:
                                  \sdramDataMasks$next  = targetMask;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$2040 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* src = "sdram_controller.py:918" *)
                      casez (\$2042 )
                        /* src = "sdram_controller.py:918" */
                        1'h1:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$2048 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                  (* src = "sdram_controller.py:620" *)
                                  casez (\$2050 )
                                    /* src = "sdram_controller.py:620" */
                                    1'h1:
                                        \sdramDataMasks$next  = 4'hf;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:973" *)
                casez (\$2052 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$2054 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                          begin
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:399" *)
                            casez (\$2060 )
                              /* src = "sdram_controller.py:399" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:402" */
                              default:
                                  (* src = "sdram_controller.py:406" *)
                                  casez (\$2062 )
                                    /* src = "sdram_controller.py:406" */
                                    1'h1:
                                        \sdramDataMasks$next  = targetMask;
                                  endcase
                            endcase
                            (* src = "sdram_controller.py:1010" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1010" */
                              1'h1:
                                  \sdramDataMasks$next  = targetMask;
                            endcase
                          end
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$2064 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$2066 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* full_case = 32'd1 *)
                            (* src = "sdram_controller.py:613" *)
                            casez (\$2072 )
                              /* src = "sdram_controller.py:613" */
                              1'h1:
                                  /* empty */;
                              /* src = "sdram_controller.py:616" */
                              default:
                                  (* src = "sdram_controller.py:620" *)
                                  casez (\$2074 )
                                    /* src = "sdram_controller.py:620" */
                                    1'h1:
                                        \sdramDataMasks$next  = 4'hf;
                                  endcase
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramDataMasks$next  = 4'hf;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \pageColumnIndex$next  = pageColumnIndex;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:853" *)
                casez (\$2076 )
                  /* src = "sdram_controller.py:853" */
                  1'h1:
                      (* src = "sdram_controller.py:855" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:855" */
                        1'h1:
                            \pageColumnIndex$next  = targetColumnAddress;
                      endcase
                endcase
                (* src = "sdram_controller.py:872" *)
                casez (\$2078 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:913" *)
                      casez (\$2080 )
                        /* src = "sdram_controller.py:913" */
                        1'h1:
                            \pageColumnIndex$next  = \$2083 [7:0];
                        /* src = "sdram_controller.py:915" */
                        default:
                            \pageColumnIndex$next  = 8'h00;
                      endcase
                endcase
              end
          endcase
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:973" *)
                casez (\$2085 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$2087 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* src = "sdram_controller.py:1010" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1010" */
                              1'h1:
                                  \pageColumnIndex$next  = targetColumnAddress;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$2089 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$2091 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            \pageColumnIndex$next  = \$2094 [7:0];
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \pageColumnIndex$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlRdIncAddress$next  = ctrlRdIncAddress;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:872" *)
                casez (\$2096 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      \ctrlRdIncAddress$next  = 1'h1;
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$2098 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      \ctrlRdIncAddress$next  = 1'h0;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlRdIncAddress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:669" *)
    casez (targetBankAddress)
      2'h0:
          \targetBankCanPreCharge$next  = bankController0_bankCanPreCharge;
      2'h1:
          \targetBankCanPreCharge$next  = bankController1_bankCanPreCharge;
      2'h2:
          \targetBankCanPreCharge$next  = bankController2_bankCanPreCharge;
      2'h?:
          \targetBankCanPreCharge$next  = bankController3_bankCanPreCharge;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \targetBankCanPreCharge$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    ctrlRdDataOut = 24'h000000;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:814" *)
          casez (errorState)
            /* src = "sdram_controller.py:814" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:817" */
            default:
              begin
                (* src = "sdram_controller.py:872" *)
                casez (\$2100 )
                  /* src = "sdram_controller.py:872" */
                  1'h1:
                      ctrlRdDataOut = sdramDqOut[23:0];
                endcase
                (* src = "sdram_controller.py:920" *)
                casez (\$2102 )
                  /* src = "sdram_controller.py:920" */
                  1'h1:
                      ctrlRdDataOut = sdramDqOut[23:0];
                endcase
              end
          endcase
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlWrIncAddress$next  = ctrlWrIncAddress;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:967" *)
                casez (\$2104 )
                  /* src = "sdram_controller.py:967" */
                  1'h1:
                      (* src = "sdram_controller.py:969" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:969" */
                        1'h1:
                            \ctrlWrIncAddress$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$2106 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* src = "sdram_controller.py:1063" *)
                      casez (\$2108 )
                        /* src = "sdram_controller.py:1063" */
                        1'h1:
                            \ctrlWrIncAddress$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlWrIncAddress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramDqWRn$next  = sdramDqWRn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:973" *)
                casez (\$2110 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$2112 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            \sdramDqWRn$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$2114 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$2116 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            \sdramDqWRn$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramDqWRn$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \sdramDqIn$next  = sdramDqIn;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:973" *)
                casez (\$2118 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$2120 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            \sdramDqIn$next [23:0] = ctrlWrDataIn;
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$2122 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      \sdramDqIn$next  = \$2124 ;
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \sdramDqIn$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \ctrlWrInProgress$next  = ctrlWrInProgress;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:950" *)
          casez (errorState)
            /* src = "sdram_controller.py:950" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:953" */
            default:
              begin
                (* src = "sdram_controller.py:973" *)
                casez (\$2126 )
                  /* src = "sdram_controller.py:973" */
                  1'h1:
                      (* src = "sdram_controller.py:1002" *)
                      casez (\$2128 )
                        /* src = "sdram_controller.py:1002" */
                        1'h1:
                            (* src = "sdram_controller.py:1010" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1010" */
                              1'h1:
                                  \ctrlWrInProgress$next  = 1'h1;
                            endcase
                      endcase
                endcase
                (* src = "sdram_controller.py:1015" *)
                casez (\$2130 )
                  /* src = "sdram_controller.py:1015" */
                  1'h1:
                      (* full_case = 32'd1 *)
                      (* src = "sdram_controller.py:1054" *)
                      casez (\$2132 )
                        /* src = "sdram_controller.py:1054" */
                        1'h1:
                            /* empty */;
                        /* src = "sdram_controller.py:1056" */
                        default:
                            (* src = "sdram_controller.py:1059" *)
                            casez (cmdCompleted)
                              /* src = "sdram_controller.py:1059" */
                              1'h1:
                                  \ctrlWrInProgress$next  = 1'h0;
                            endcase
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \ctrlWrInProgress$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    \refreshCmdIndex$next  = refreshCmdIndex;
    (* src = "sdram_controller.py:708" *)
    casez (sdramCtrlr_state)
      /* \amaranth.decoding  = "InitOp/0" */
      /* src = "sdram_controller.py:709" */
      3'h0:
          /* empty */;
      /* \amaranth.decoding  = "ConfigurationOp/2" */
      /* src = "sdram_controller.py:734" */
      3'h2:
          /* empty */;
      /* \amaranth.decoding  = "Idle/3" */
      /* src = "sdram_controller.py:784" */
      3'h3:
          /* empty */;
      /* \amaranth.decoding  = "ReadOp/5" */
      /* src = "sdram_controller.py:809" */
      3'h5:
          /* empty */;
      /* \amaranth.decoding  = "WriteBurstOp/6" */
      /* src = "sdram_controller.py:944" */
      3'h6:
          /* empty */;
      /* \amaranth.decoding  = "RefreshOp/4" */
      /* src = "sdram_controller.py:1089" */
      3'h4:
          (* full_case = 32'd1 *)
          (* src = "sdram_controller.py:1092" *)
          casez (errorState)
            /* src = "sdram_controller.py:1092" */
            1'h1:
                /* empty */;
            /* src = "sdram_controller.py:1095" */
            default:
              begin
                (* src = "sdram_controller.py:1096" *)
                casez (\$2134 )
                  /* src = "sdram_controller.py:1096" */
                  1'h1:
                      (* src = "sdram_controller.py:1098" *)
                      casez (cmdCompleted)
                        /* src = "sdram_controller.py:1098" */
                        1'h1:
                            \refreshCmdIndex$next  = 1'h1;
                      endcase
                endcase
                (* src = "sdram_controller.py:1101" *)
                casez (\$2136 )
                  /* src = "sdram_controller.py:1101" */
                  1'h1:
                      (* src = "sdram_controller.py:1103" *)
                      casez ({ \$2142 , \$2138  })
                        /* src = "sdram_controller.py:1103" */
                        2'b?1:
                            /* empty */;
                        /* src = "sdram_controller.py:1105" */
                        2'b1?:
                            \refreshCmdIndex$next  = 1'h0;
                      endcase
                endcase
              end
          endcase
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \refreshCmdIndex$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    (* src = "sdram_controller.py:670" *)
    casez (targetBankAddress)
      2'h0:
          \targetBankRefreshCounter$next  = bankController0_bankREFIcyclesCounter;
      2'h1:
          \targetBankRefreshCounter$next  = bankController1_bankREFIcyclesCounter;
      2'h2:
          \targetBankRefreshCounter$next  = bankController2_bankREFIcyclesCounter;
      2'h?:
          \targetBankRefreshCounter$next  = bankController3_bankREFIcyclesCounter;
    endcase
    (* src = "/home/lpnm/Documents/Electronica/FreeFPGATools/oss-cad-suite-linux-x64-20220517/oss-cad-suite/lib/python3.8/site-packages/pyhdl/amaranth/amaranth/hdl/xfrm.py:519" *)
    casez (clkSDRAM_rst)
      1'h1:
          \targetBankRefreshCounter$next  = 10'h000;
    endcase
  end
  assign \$831  = \$832 ;
  assign \$1180  = \$1181 ;
  assign \$1193  = \$1194 ;
  assign \$1204  = \$1205 ;
  assign \$1215  = \$1216 ;
  assign \$1224  = \$1225 ;
  assign \$1235  = \$1236 ;
  assign \$1248  = \$1249 ;
  assign \$1255  = \$1256 ;
  assign \$1264  = \$1265 ;
  assign \$1279  = \$1280 ;
  assign \$2082  = \$2083 ;
  assign \$2093  = \$2094 ;
  assign clkSDRAM_clk = 1'h0;
  assign clkSDRAM_rst = 1'h0;
  assign targetMask = 4'h8;
  assign targetRowAddress = ctrlAddress[20:10];
  assign targetBankAddress = ctrlAddress[9:8];
  assign targetColumnAddress = ctrlAddress[7:0];
  assign sdramClk = 1'h0;
  assign \$33  = refreshCmdIndex;
  assign \$57  = refreshCmdIndex;
  assign \$121  = refreshCmdIndex;
  assign \$179  = refreshCmdIndex;
  assign \$205  = sdramClkEn;
  assign \$223  = sdramClkEn;
  assign \$277  = sdramClkEn;
  assign \$331  = sdramClkEn;
  assign \$333  = refreshCmdIndex;
  assign \$341  = sdramClkEn;
  assign \$347  = sdramClkEn;
  assign \$353  = sdramClkEn;
  assign \$361  = sdramClkEn;
  assign \$369  = sdramClkEn;
  assign \$375  = sdramClkEn;
  assign \$379  = sdramClkEn;
  assign \$391  = sdramClkEn;
  assign \$397  = sdramClkEn;
  assign \$413  = sdramClkEn;
  assign \$419  = sdramClkEn;
  assign \$433  = sdramClkEn;
  assign \$439  = sdramClkEn;
  assign \$445  = sdramClkEn;
  assign \$457  = sdramClkEn;
  assign \$463  = sdramClkEn;
  assign \$477  = sdramClkEn;
  assign \$485  = sdramClkEn;
  assign \$497  = sdramClkEn;
  assign \$503  = sdramClkEn;
  assign \$511  = sdramClkEn;
  assign \$517  = sdramClkEn;
  assign \$525  = sdramClkEn;
  assign \$527  = refreshCmdIndex;
  assign \$531  = sdramClkEn;
  assign \$535  = sdramClkEn;
  assign \$545  = sdramClkEn;
  assign \$559  = sdramClkEn;
  assign \$563  = sdramClkEn;
  assign \$565  = sdramClkEn;
  assign \$577  = sdramClkEn;
  assign \$581  = sdramClkEn;
  assign \$595  = sdramClkEn;
  assign \$599  = sdramClkEn;
  assign \$611  = sdramClkEn;
  assign \$615  = sdramClkEn;
  assign \$619  = sdramClkEn;
  assign \$631  = sdramClkEn;
  assign \$635  = sdramClkEn;
  assign \$647  = sdramClkEn;
  assign \$653  = sdramClkEn;
  assign \$663  = sdramClkEn;
  assign \$667  = sdramClkEn;
  assign \$673  = sdramClkEn;
  assign \$677  = sdramClkEn;
  assign \$683  = sdramClkEn;
  assign \$685  = refreshCmdIndex;
  assign \$687  = sdramClkEn;
  assign \$691  = sdramClkEn;
  assign \$695  = sdramClkEn;
  assign \$699  = sdramClkEn;
  assign \$705  = sdramClkEn;
  assign \$711  = sdramClkEn;
  assign \$715  = sdramClkEn;
  assign \$717  = sdramClkEn;
  assign \$729  = sdramClkEn;
  assign \$733  = sdramClkEn;
  assign \$747  = sdramClkEn;
  assign \$751  = sdramClkEn;
  assign \$755  = sdramClkEn;
  assign \$759  = sdramClkEn;
  assign \$771  = sdramClkEn;
  assign \$775  = sdramClkEn;
  assign \$787  = sdramClkEn;
  assign \$793  = sdramClkEn;
  assign \$797  = sdramClkEn;
  assign \$803  = sdramClkEn;
  assign \$807  = sdramClkEn;
  assign \$813  = sdramClkEn;
  assign \$815  = refreshCmdIndex;
  assign \$817  = sdramClkEn;
  assign \$914  = sdramClkEn;
  assign \$920  = sdramClkEn;
  assign \$926  = sdramClkEn;
  assign \$928  = sdramClkEn;
  assign \$940  = sdramClkEn;
  assign \$954  = sdramClkEn;
  assign \$958  = sdramClkEn;
  assign \$970  = sdramClkEn;
  assign \$982  = sdramClkEn;
  assign \$988  = sdramClkEn;
  assign \$994  = sdramClkEn;
  assign \$1000  = sdramClkEn;
  assign \$1006  = sdramClkEn;
  assign \$1012  = sdramClkEn;
  assign \$1014  = sdramClkEn;
  assign \$1026  = sdramClkEn;
  assign \$1040  = sdramClkEn;
  assign \$1044  = sdramClkEn;
  assign \$1056  = sdramClkEn;
  assign \$1068  = sdramClkEn;
  assign \$1074  = sdramClkEn;
  assign \$1080  = sdramClkEn;
  assign \$1086  = sdramClkEn;
  assign \$1092  = sdramClkEn;
  assign \$1098  = sdramClkEn;
  assign \$1100  = sdramClkEn;
  assign \$1112  = sdramClkEn;
  assign \$1126  = sdramClkEn;
  assign \$1130  = sdramClkEn;
  assign \$1142  = sdramClkEn;
  assign \$1154  = sdramClkEn;
  assign \$1160  = sdramClkEn;
  assign \$1166  = sdramClkEn;
  assign \$1174  = sdramClkEn;
  assign \$1187  = sdramClkEn;
  assign \$1271  = refreshCmdIndex;
  assign \$1284  = sdramClkEn;
  assign \$1300  = sdramClkEn;
  assign \$1314  = sdramClkEn;
  assign \$1318  = sdramClkEn;
  assign \$1330  = sdramClkEn;
  assign \$1342  = sdramClkEn;
  assign \$1348  = sdramClkEn;
  assign \$1352  = sdramClkEn;
  assign \$1358  = sdramClkEn;
  assign \$1372  = sdramClkEn;
  assign \$1378  = sdramClkEn;
  assign \$1392  = sdramClkEn;
  assign \$1400  = sdramClkEn;
  assign \$1408  = sdramClkEn;
  assign \$1410  = refreshCmdIndex;
  assign \$1420  = sdramClkEn;
  assign \$1426  = sdramClkEn;
  assign \$1440  = sdramClkEn;
  assign \$1446  = sdramClkEn;
  assign \$1460  = sdramClkEn;
  assign \$1468  = sdramClkEn;
  assign \$1476  = sdramClkEn;
  assign \$1478  = refreshCmdIndex;
  assign \$1488  = sdramClkEn;
  assign \$1494  = sdramClkEn;
  assign \$1508  = sdramClkEn;
  assign \$1514  = sdramClkEn;
  assign \$1528  = sdramClkEn;
  assign \$1536  = sdramClkEn;
  assign \$1544  = sdramClkEn;
  assign \$1546  = refreshCmdIndex;
  assign \$1556  = sdramClkEn;
  assign \$1562  = sdramClkEn;
  assign \$1576  = sdramClkEn;
  assign \$1582  = sdramClkEn;
  assign \$1596  = sdramClkEn;
  assign \$1604  = sdramClkEn;
  assign \$1612  = sdramClkEn;
  assign \$1614  = refreshCmdIndex;
  assign \$1640  = sdramClkEn;
  assign \$1674  = sdramClkEn;
  assign \$1714  = sdramClkEn;
  assign \$1728  = sdramClkEn;
  assign \$1740  = sdramClkEn;
  assign \$1752  = sdramClkEn;
  assign \$1774  = { 1'h0, \$1772  };
  assign \$1786  = { 1'h0, \$1784  };
  assign \$1794  = refreshCmdIndex;
  assign \$1812  = sdramClkEn;
  assign \$1826  = sdramClkEn;
  assign \$1840  = sdramClkEn;
  assign \$1854  = sdramClkEn;
  assign \$1868  = sdramClkEn;
  assign \$1882  = sdramClkEn;
  assign \$1896  = sdramClkEn;
  assign \$1910  = sdramClkEn;
  assign \$1924  = sdramClkEn;
  assign \$1938  = sdramClkEn;
  assign \$1952  = sdramClkEn;
  assign \$1966  = sdramClkEn;
  assign \$1980  = sdramClkEn;
  assign \$1994  = sdramClkEn;
  assign \$2008  = sdramClkEn;
  assign \$2022  = sdramClkEn;
  assign \$2050  = sdramClkEn;
  assign \$2062  = sdramClkEn;
  assign \$2074  = sdramClkEn;
  assign \$2136  = refreshCmdIndex;
endmodule

(* \amaranth.hierarchy  = "top" *)
(* top =  1  *)
(* generator = "Amaranth" *)
module top(sdramClkEn, sdramRASn, sdramCASn, sdramWEn, sdramCSn, sdramAddress, sdramBank, sdramDqOut, sdramDqIn, sdramDqWRn, sdramDataMasks, ctrlReady, ctrlWrAddress, ctrlWr, ctrlWrDataIn, ctrlWrIncAddress, ctrlRdAddress, ctrlRd, ctrlRdDataOut, ctrlRdIncAddress, sdramClk
);
  (* src = "sdram_controller.py:222" *)
  input ctrlRd;
  wire ctrlRd;
  (* src = "sdram_controller.py:221" *)
  input [20:0] ctrlRdAddress;
  wire [20:0] ctrlRdAddress;
  (* src = "sdram_controller.py:223" *)
  output [23:0] ctrlRdDataOut;
  wire [23:0] ctrlRdDataOut;
  (* src = "sdram_controller.py:224" *)
  output ctrlRdIncAddress;
  wire ctrlRdIncAddress;
  (* src = "sdram_controller.py:213" *)
  output ctrlReady;
  wire ctrlReady;
  (* src = "sdram_controller.py:216" *)
  input ctrlWr;
  wire ctrlWr;
  (* src = "sdram_controller.py:215" *)
  input [20:0] ctrlWrAddress;
  wire [20:0] ctrlWrAddress;
  (* src = "sdram_controller.py:217" *)
  input [23:0] ctrlWrDataIn;
  wire [23:0] ctrlWrDataIn;
  (* src = "sdram_controller.py:218" *)
  output ctrlWrIncAddress;
  wire ctrlWrIncAddress;
  (* src = "sdram_controller.py:205" *)
  output [10:0] sdramAddress;
  wire [10:0] sdramAddress;
  (* src = "sdram_controller.py:206" *)
  output [1:0] sdramBank;
  wire [1:0] sdramBank;
  (* src = "sdram_controller.py:202" *)
  output sdramCASn;
  wire sdramCASn;
  (* src = "sdram_controller.py:204" *)
  output sdramCSn;
  wire sdramCSn;
  (* src = "sdram_controller.py:199" *)
  output sdramClk;
  wire sdramClk;
  (* src = "sdram_controller.py:200" *)
  output sdramClkEn;
  wire sdramClkEn;
  (* src = "sdram_controller.py:210" *)
  output [3:0] sdramDataMasks;
  wire [3:0] sdramDataMasks;
  (* src = "sdram_controller.py:208" *)
  output [31:0] sdramDqIn;
  wire [31:0] sdramDqIn;
  (* src = "sdram_controller.py:207" *)
  input [31:0] sdramDqOut;
  wire [31:0] sdramDqOut;
  (* src = "sdram_controller.py:209" *)
  output sdramDqWRn;
  wire sdramDqWRn;
  (* src = "sdram_controller.py:201" *)
  output sdramRASn;
  wire sdramRASn;
  (* src = "sdram_controller.py:203" *)
  output sdramWEn;
  wire sdramWEn;
  sdramController sdramController (
    .ctrlRd(ctrlRd),
    .ctrlRdAddress(ctrlRdAddress),
    .ctrlRdDataOut(ctrlRdDataOut),
    .ctrlRdIncAddress(ctrlRdIncAddress),
    .ctrlReady(ctrlReady),
    .ctrlWr(ctrlWr),
    .ctrlWrAddress(ctrlWrAddress),
    .ctrlWrDataIn(ctrlWrDataIn),
    .ctrlWrIncAddress(ctrlWrIncAddress),
    .sdramAddress(sdramAddress),
    .sdramBank(sdramBank),
    .sdramCASn(sdramCASn),
    .sdramCSn(sdramCSn),
    .sdramClk(sdramClk),
    .sdramClkEn(sdramClkEn),
    .sdramDataMasks(sdramDataMasks),
    .sdramDqIn(sdramDqIn),
    .sdramDqOut(sdramDqOut),
    .sdramDqWRn(sdramDqWRn),
    .sdramRASn(sdramRASn),
    .sdramWEn(sdramWEn)
  );
endmodule

